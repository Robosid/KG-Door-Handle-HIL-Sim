// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gSQzccQCfL2Nnn4WVVTKBYR98OfvTXrksz1QvxcLJ3linwNbZmflQ+v/ovFWV3hiGMmIhco2x13A
NPaNCrpIvMhX0pIOrK/ChkxJL0uVKIi3aKMMNgdoLxV1hVWDdPm5mLyR5XbaEgQN0JQ2H/WsIkF+
hlmSpgj3qJFKhW4hoVm+AHRF+AUGV7e/HOCB61J3JI6FeR2zyGfSBeBHEUnCNBVvlO+Xe3TShDK5
PnaOHB5Kq4D/C35lTdsnuoH/BMFAwSHjpK+lnUKpi9FdagGSclM6kTi4cQyeKt8OabINIHDjOjSI
Vv+o2nPOsOM+2tAQT3z51MmG/lvkjmyBnTVy6A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6368)
xm5pD2twh+aD2fGBbe0qsOu5I2gPVPPgZOZ1khrNakEW+L0xQcNbt6qUsozZdp+6VDwo1ILDIHgs
/Klftk04WhjmMWxZlAkPf/Qie+QbFbPQrv/g5lHmfkVjMV55J+QBfO9Z4+kFvk73L7CAel3W8g9c
HkI/QWn35P5g/AyRlPcyDcvje4x01LpQg7o3WodQjtdKsO5xV0LBa8aBep3rfQ9Arn4DQLiWTP7c
Rysvw5EpMjXPsa3zn0UDN5DJHejqFJeap4FkFL1NOEaY46RzFDatLAU0hzCQuajrT4SgLQUk5/Es
AzbfTY2czHpKKGCmCqkzBP2E9VUaN2xvvT95wazDS2v23XbJL7lc/IAG3C4BY6R5rqsm5JBU8BOk
0P1exRMTbV/nbpjPl9sgVJE9jzrzancI7uwrT1eZwpktt9YO4fDHSiOMq3ykLduD9iybM5hbTQWn
o24XJZW7ltFC2iWU86Unva9lE7R5/i2OmbDhjP2CRA0TKMJsq1C1n2Ah+fINvGZesB7xR551OfIO
CjcubmmHi6BULY00G3aKFoNbLxW1YvMuljqDvGzz4gzyy7mBhFHdNy1PX4IOyPV4BTNYCB7o0yJu
brhtXgyMi7nvhJy80G/LOTtcF9/xMj2a/PzkDhRTT8UmicV3NgxB3vOtV5GV6cQXnlBYjiRXYxm2
VsjdDbngVOuO2BwLTduNpf+6a2hnO6ye2SHNOH6DToPnLc2EBHsiD0R9SC/WM/WjJ3E+5N1ZIOTJ
tfG7u7Q8It1Pu3sMvAhYAfhQm2g7jtjZZxwUxCc4lL+147kBjWnmFabynhRHMp46blIvIvjEldgv
EYnft+zYaP7jE9Py1B7YDqN7SQ9IH26kDnXmt/YjBSEB5VzqUpKto5JgVFpOibJa8ZcrRcl9iA90
IIOvIz6nwuUjRFlcInvfmy+63n1cssG4XnlayXiICggZhat/aUXZbZs9Pu5VayWWBQiTiWFSHGVe
unT1CfFMhN0piE6ljfhsR4UsPvcjMcq7CszqfNBF4hFvbmxzIWd4EqxqrF0AXaLbLBhRt+r1UJ7h
CjAAOuLLziQoeKp6nBQsDZQqNQBJqeSOMOLbySp8EPOD6c5rml4zc/P69DayjpP/lvI52o1ITNLI
d3bYKSuckXKtH8AWxz0iG1csLYcf3k1ks+5sPRnyA9BpeTIDh7B6I8qqldGaw+uY1+yqb6M8PEQn
NTMUKzP/hQtPk+tkfgpDjExqC58lg29EOYeNb9dxrT8dYGgK6mE3G30QhVQXJKZqznH6xdx+/it7
o5Lw/xh4ajkjT72SQAQ0s6jb5vgZsd9dUS+diLEJFszsZ1vj6HZUTlxeWVJi5F0KwcfeTGR59hbt
9OcyGT765nyUJfqe+JbL7u2RdJ2mg75TxjPYrcgjaVOUotkVWxa31dOftD2IOCYTJQ8RhzUvkyC9
IW/ul5wfpTkjPNFm/C4fJ0MGf82XmHEtbhBeIU9fqFjT07y36IrI+ErcyvTJzUm2mrHLe/Uxn+B4
urpTKF77YEI06mmTAqQrqIBAJH4VuOMMWLfIWFjDpPUlFL8UvydPO9dkN8CIhiam4TRyMYADSI0N
je68wo2ynLGAVpzxVVwaeVTGqr/Ex6EwhIIr5Q6mTDPtDqrFoZL/lGb6tjjIaG27XLIGG11sZ8rS
eMy11E5nr59HRpbfz5BJ4UauxDULiKI5n9QPG8ofxGo64xkbGThZoRevPY90qQbe9DKdgLRFRjos
U9sgHMyV5XZv9fAC6ZYdEpcbwAYX9R1SaGHdf49pZNDbE9VHP9WMOnuYZLWq9gvZ5qKUOba5oSwg
bTod7HLKRubMoDeuC71qapFeOEb/rE2wQJnyISpBU+EMp4ZYAHIVtxsMlAb7cAKljMq1AZJaumAO
5fpYgwtC9Te2r7yR26h4te+OAenRw6jFCKRkw2lNwQvhI4vLVovhuVJNG4acdwsMX6HuIzkGvj38
XGYhQLDuoK2vhEhNqR6UX0a3FnliFjJNq9RdK0N9V02Czd0nKvU7cxw1HwlUIkXzaWtfGnVC2yym
OFhtKVCgf3MN7x3MuvsrOLsblaXZrj+ro9HZB8gHwQ737jFM5BdHQBAVj8ad4tLfYN/IDkwQHkbF
848gGSSrC9iuquEhH1/XvtPONQkEI98K9GlZ1eUb3uv31Mf7L9fj9+5gl88BpraaRlm43Mf40Dr/
0Y12ngYlHExKaZtldTbYZ7tceNg0WoZDZY6+Wr/Yk0R5zPDIBgcVJgk6rBAb+aOjw7OhX1hZtwXQ
b6lgjv+kQ/phzjpS/DtMw7605XWUfwckrq7Y02gqVInHplyJNZ/tsMHWNtWKTArd9D8vuzh+4rGr
UzZ/kRz7P6RWFBQLPoq8CdabRfYaDXp2m5+DmOcDZ7T28fhKuGtlM0bZ9mcuB3FutE3Gb0yFQsYK
Kigm78Hcb39goZIYzP1yqJqyYV7PUMae5Kon4u2WN5jHJX9V6qqYhv/NBTI+XPsZ8kc8kpNp8fxa
x4RSFJf709gBGReaPxVhrKtFdf72oEDJPMPCoQXAPhH+Yvzgovo1S+WdZ4oCQIpL0SPJzDWrYAk6
4NvlU66DdNnqf+PpODkzOnfLt3dDptCtG+zSNjAVc9KWmMj9+8gz5Kocq8HFEVW88ecVwhTfIAyG
LtDVAJDgj+WQF29YwnQJPKhNPOfR+3LQ8pGIeRzAikP9kXv1viobnlPZ/cGgN2MfZTmdO40iKsXo
xEQxcI28NuVc8e+Yq7WysdqYWPzwESidaPnqq4pyG238S8Eodhd3QxhzW4Mp9+YBxAq/ietUpwzc
UI//7ucPLQqP8ijeDyNSMxEjXXxzU2jyazqqVjMDsrGFCzKlLeewsfODwshptqvcnkKPRl7mHs7m
vbYgzjARulC/NIlk0rgxupRUmmU/gJEXAvVX3av30S6teC/8UmyB8YTqvQUNP4loZvtHppVDhRSx
+qCi3ZWPZ2815Be8mOGs6s+rgkd9erbYmtVVGywudBVT6UwMp2cOpuwXtG56JWbr/I6QArmCR/MA
53c5ERpPrMsA38y89GDFZLYm1uLQMU+WNYPzJeJm3gYlixBC4ZEawTziOx3kIAp2IVIt/TqCOG0B
KR5jpII4GWHMU76BJyToqk6Xr6/cAnBAR0gxCH/8PyL8dHhZ7KBgpk7yEeiThr6ydPWzWTnXZt9f
hLQDtghwTiOwEd3Y537tmUc1vQ9A/LjMZDVHFI5XIwkaWS1QU9DHj19PiX/cx+EregRAiaUaKiI+
FDeh1Q/2JPb7CUCzYcbsbvPlpmEWt1WOqMict3xxUULvxAqZfUBjB3aWn785173dDXn8L5DjI7zY
kwDAdS8pMsNMaYD376R0+8dknE2bUpQwhdo2/jdXlEoulRBeC392JAWwmnK+Q4eqSHw/xiZ0J22o
Y198UbJtIwuge2aV0ZzCs5NcKGHNJ3pIXQSAXb8lV65MFuE4NRZtR7DjzL4X46aAPstSfil3ji4O
ihZlf9QS5fHPvztBHLBqfGKPk+9F11sD1FsvhgjzTDm8aWlDEJRdihwOAZC2V8RH5ntY1vnKFWxW
dd+E8an3XzOtpTfw8RL6LbJm6U3OpzEN2h3O9TtIWFSOPz7y9Fm9FgX4D13cR+OQQDQVXEf4gIpO
jF9bO6buxg828cizKKD/RzzL+PbVfquOhR/lRw4flWKE+IoD5Aes9paJfmTQaZkpCWlDsNYkClEo
lqh3e7DDHQCIP9oNqzVknlV9Z5VgGsOXe15CADkd2Y3MYx9M20i7dLv82eUdIByAFVXCHr9/HnKh
O73EZ1VdYk7ca1TsdFYd9GkN5ZKS+tY5IPoH+M2KZEHDmvzIRb3H6/XkdXj/HjbsxN1pnhpmZEpy
95pI6Rz5vhuQu6sYQIW3q/1FrKxa4OP+r4UnIV9NHzZLDP3wkanQw+YLBzZ4wCvlVFR0uijEHuUJ
o95v6LJe1q3HeqTP+xKeWffUJ0wMzbPbPQCpIJ4rJJJ+/P8fwG83KM9ir2q3aPa3gHOC8/IioK5H
uRueeTqtp64AlNyxqO2ckaVa+3BGgM/DBhNiA+BqQ+KgXBXBs9R0icjzuVpOivpkuXIq9bexaatm
c6uIQ+TBrrRnoUTfGAeAuORFvWYoXhhfXNf/s/cWDPsToemvKFIytSmKVbVNXDiR/KHyQEidHd46
WyilR7M1R7b31OgdGmAlMx84YxKXn6b/pvaINk8payvHqaeyVo+g3ZX4Cg3jRzAnG5bExuvvGGOv
DGOuUfK9USsl4hi/CvEQh1gHcByt96yVE5dy9UoGNAjDzVJBxfIf0q6PcWg/tWrIFe6ptyo7QgSJ
8QFBT3mLIRqjyZC8rCS08bxO3+6zMVglBP0rHZ0wOB9P7UenS2+G1nUxbtgMgUdX55g2nfY9zIuw
Ue7+kN9BHr/wu66tjTzJunVVK6jFKfrmaSBX7HOz6Zd/gXK3Q0KFgIGs+3NASP6uIHAL6RC14a4L
KjOPukTAdwp2haHTZFOPBHhYdR5ref7UylZyRhY3R1kFb7uXJ71MsdzZEy08iUsGF7PNlndkDBtm
IRZ2WH7JoD6p84N30IUFKG9IntSwLQZ8+HjcXdQlpoqKMeFUMobXcH4ELW/4TU+zriwC1T1N8mBQ
P7WGdOUPsM747ZLZfjtpC2EB4p/OmB1eev5EOfd/d2dQBcaT+qzG5KiDV/BkmC2i2DHkKjN535Ar
n6kW1a/a2QVRiofZXofUADWKg60tYJcTlReDKcPwzaWROYcsu9t0dsJd3zUgEl9eta84LY4m8eri
2JlomWwvemJcfISyc1BQBBR/1fNMxe3m36hnhsDMy1yXRC4Ft/Jly4MOABJtA+6mrS30ybLEUkvg
wDgZpn9h3Ct2xzu5ZpKvfNxtTCHecJHDf6WkE/hoeKxc0rCq5ATfONi4fOp7w1qtEHyd3XH4CBtd
QGqEYMRoEw1ctISIx2yoyzD5OODcQEDcls74q7F+Us38WSBJwi8gCh2LRSZ4FGD6SgwAZP6kIoDm
Hh8XbIz1Rv+9uHf9iEClAI2xR3aaHFVC1+FgK6qVzpOMB+L3fhPAVPX4ouUS8tAPBXq/vtsprX3b
uBCnlbMDIgC3D6H+iFgcoUf3C/b7Lf5ATekWQa9hw+cbU2LHcz125sQqAApx3F1apNK1T4xfvOOj
83ZTgDQVKTruBmh1XpNdiiFs4Wlu07jvBewXiU5rgb+/kb9R+T5cGwp1TzxKh/c0WEDBjGcGbuCu
1ny78Qus5e/qR2Cq7Q+z1hzvmI3BXIC/0LA5Uz987AWvU4epPEk+VmLvzOSxyrb99Z+t3TRoMzth
5/amQxEAWbHd0m7u7uFxAreypbywSNDg1iZj+T9SGcWJCNKrEolxLlDCTT5BOtKttZnNnKDrPpdS
tLiP8vH3ZJusq/XrjKUS0DIgdccqrxvLv7qMzpuUc5Oft0hzAQUsadZ/0rySc7kLUaxEE9AXQ0Hy
CWv10iFWUN3W3cZJk0SF1FnFmDFKmQEWpsLQxEkUKZtY3Zwq3aUZOCBpGGt1+Os5KoFo7dhTkkES
F18pJgK2CbdbXOAogIRKQX9fT+KRTHdqRtqPE6xFJzlBMArYfYNZwe3aKkFsEsTkncqGl9GWVIT1
I9t83gUajwKq1Mw+GLss60mDGiEBbWXJLcktc0CzvwpU9ynPdrRZDxKOH3KCmuaHHYTmwfi1kKTw
K54SeTU+i2WqoVFu90GX5Ct8HxRZMIO4hG5+ZgxUO4xSDVWCdBWHE9rndqXJGDY57Jltcql1feOq
RMXZElIoJjY/8ySK6ReBLAABNKRL8PM51jjdvG5huRKYmIaE0K52k8TNb8eyEjlwyp4O2jmRIdGs
L3qroYgGqu05bQyGitqcC3NSUhGrfoIPpkd4pliC+ghOzILDOIJdvv7PCSbItxujFFJHBVmjbiRW
68q/r/NmBCA0WT1kL5SA/t1z/v6t6IbiB+mBqMLg8hwUyNTJSJ0gdnmFEPImZSuTH2sRZ4F5mLyz
EteRcm9fUoDt+fBW5UEhHeBpY10K5UYAmqrNE8aSPnxVPzGu3wzatdpf384cfsJJLxm0Qb9vXxP+
o4jcxucmfFQ0bJvIiLj+LyCx80ijj0lGvlZLiPx0oaTAxqTcUjhJI42DOdXDaXvr7B8ll2mvxOb8
uLC4OUoiP50yDN1VQ1hjDvi+VjjfQfPj11Df8kasOhmDMPqBVlKCLuZCcjqZE2QVuSd/bGrRsEW0
uc9w+DH1Y9f1TDzxAIZjQ/vAc1y0G6zr2lV2a55ncA9stXKiC1QdGg424N9fc43ZWnoGgY8x6JoM
do98/Wie099AQs9hUVyUtrhDq60VWACjUFKkPWPWrVR3+CTxeSjvwh/J9RA4IQu5fIjzG4iCfj0G
ZQ+SniblzAa1oVlIVSf5fJy0R6uf08Tm0pOHPJOTJ7b6v+QPMknfWzq6zVQxpnDUa847QDbMT5Kp
cWVxrdq4qPve3S2uA3B4NnVqoiFtAbgK4ebnDbpsD6Ntldp56wIrJqOKhrmgeWfgvEF2zh9JmQJR
BtJ5i9ea4dRgVwLNWb7MGchnQy7KNMojRPlsbgslQj13VWfNRZZC0SstgdOlho5Fbnk2KL6CkQxk
BG1Gc1wKscbX53MzK8zX1F+blSc6DODrb6ZP6c1FqKqfm1qNAIV3wz3Y29MLQSCU2Hf0xn38vabM
6AM68whDA7P9zqbWHm63mnOdINf9r6FQ/D/xZhn47p2HXRBzjXSKuqRM2zWOviS7fHJXiQFMyK9G
XkZnDE+rZUOIqtIDTaRPZSUw4WxuT3jNiXGysAysSBTVep80Uyf4txcyQCHr/GaBBA+NPDhquN31
/WvdCkRRGSe3COMsbgUB/khmq8JgviZyYJ8mIR5uOVNTa/wuOkU96LkdYDwr4Ske04UZBM1rRDuO
lpM/yO9K1wE0diGK1QA9g3Y1F4MeU5fHvhAPvSe0ADvAiidCxaQ4bkoV8Tc1PhXKJsLBsaEdt8E/
6Nm+dcrB/oOlC1lWKm28mi8jAn5s8+6H5u1EEAd9NpHagCUnmei5SXPDr73MyA5n4koEui3ePWXT
Zxhu8s3xtrsCgcXoUCYWOmwprc+5uZhCgHh+LPtSZwKO/2XJgSXV6AGX5JnaVex3rr3X9aivEK9n
7TBg/DDClWi9uvuot3KHwQveVDX8ImS+EqHE+PNkvDmy0HghzisXi6vS8LioQdy7JOIgU7GY+SH0
iY9GxT6MzhY8/utAOSQ9zGFuEX3XSMxleSD5pXH1YuBb1vHq8pKDDpJhZH+pg68UmpACZN/9YiHk
xEPgWGTPnWYzqu5TkBlG4uu+uSZmiCRV3JqBqmz60j0ZKBXvfzNJhsq/lUbCd7hWcFxiz9pBGUZP
abt68HSdwv9ouPCFGrvVSxWkwmLZgA+TGBFcWwmKfsmKPw72V0WrWKumKW0H9bXCXAJPvOlBxUco
u/qZSy7AA/d5s/FgIPs8mrIjrVskX03/yY6jDalymg+pt20LErl9/0JQp4BYHCEuEph50sEcxnxr
PYTnDWVocTXDG7UvApk2KkW/9fHPkGwIxlLOafGEyFGJHpJdMQgwCgCf+55gzHrpNEF28wJH4tPy
BtWQgSvc7aMEd4eBqCHvlIsjEDYJLiLJbe8RtvAYGyx4OgQTVYPNzzLfoVN2Lor5FsqpFZG5nP0D
1SnSw3iEozVbToFO4ykOcDEAMoFPg0IRF4B6fGvZK1z4R3q4Eg67L1tzAeJMy8BViPCKlsgPo5mt
4y8hHHz+I/s1rtpdaecY9/QvV14B2qeVvfnF+ORP2tlBRsYNmB5R00HAPrczQuJBUyAO2wi/FPhk
WvV4ryZuQaeEoEygbZt4jsoAEFkgQISntfHlyb9LSXjx7FH4T2VcyzJLOkGc4XifjOMUK4Isx0K1
d0ZFxgqGfYHoQa+VAghBOgcLgdvLkrLUKsy1nwgYhI0GSaIX5AE1Dnximy+AkwA63hfxcbbpxBXu
xbe3U6gQK5SWWpatuh/fpha6rw3OuSYCpgFLuXHtCnxwcPiSewLCkI8tWdd1VlJXAUIz4EBm1PSf
k1bSTpQg3RY1hbKasDx2T4N/bRnXQ1ZSJD+apUlj3Cx8+iSTQlk+KPJLTMgC8Diu0bvLWPq/3ZNP
ghbt6q/MwztwRwkJP1jiEU+MhBX2BRsLrVjJeqWTYKJIYvy0lrOYvEMmM4Dc7i6zEYNOY8dj0Oaj
+pcRJ4j2Rfjjty0j0DfykK5KQCiZppkwx/c693+27kRwS++MKrLsnqHrSzVq7uyOIX/d/J5hGAGD
8cmvxom9eliLe0j6c1Z1xmuyrznNlLpPtu0wNrhxLpxIAmfBVV/TgaM4vRInZk++EiX3X9mGzZUw
LIHeLgcabmPNi5RGw8MDDM0+SdqchqaKoTbz7Zoqm4XjKXi0ggAvUQQEdan+nW3IpNY/WgfIIZvP
qi75HJ3aYK/6Q2FnIgk7y8v0uU6rWpdFopEtS/Nm2R0wdPUYN3hLWzk=
`pragma protect end_protected

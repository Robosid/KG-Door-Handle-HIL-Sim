��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��� o�tL��nàZ�m�E*��ZQW��v�#�ͻ��n� T46��н����w�89�#�u��tJ.���Q�9���q�X��Z�(��������������Η������n���j)E�i�P�\Gj�f�Dκ�9�d��k.��-�s�+F`�9r?�4L�a�l�&�o�tƨoz�<��T����[����w���}�M�r�{���GH�����Σ��	��%�� ,a�Ew���m���8�n�7�Kr��V�I�>0ڦ<��̇���v9�_�M���}	��!r��څUѤ�<&kW���q�D�\d�+yg��32D�w�^��8��A���5�q�����e'yX�N�/T]��ن�O?�䩇h��"٭�V_q��m�ʻ-�LR�����y��ϡ#�Қ���9������M��SS�
����rO$&�^�T��AVV:�N�Ԧ��儥5s�ph����&�,� �U�}���s+i� �ҝ����'ƀ�lp�� .��&���M�r�0\R"̢���Aqb.N}.>�$Z��'͎� �UP=}q�p�����sKF��y^r
W+�;�J�ǯiz�������
�ӰS�ݚ9��0��;����E�UL?��M�C��dw��8H�M��l�r}�G]P�g>K:^a/[��h#��k�:�������T:�y�.�v���z�C�J�]M"K�*Z_����}��wm���jk���6y����F�u/��-Y��ޓ���_���`/x���%�u8'=��фԒ
��F��^|�z��X��������rw�z�{
5��w�_st��x�$}�f�#D���+��E��[�׌c%~=E���Gʡ+�2�� ��I�.��j}�!���O;��s˟��k�p^��`"��hU݆�-�@"B��#�z��:�
�|�j�*)���4i&\��9��:�yb2	��NT�b"�U�<�K�9\`�X��-_�Aj���:lSt$6���1��ol��=S�Z�Z�ψ;3}Z��e��̐ˬԖQN���-ߧ	H�$�f)�@u>n�ny���{}<f|#@@�e��q-n.���얛��]�g%�ȍ}Lg�0�֪���]q�O��\�'Ln�(C���x���i�8Q�u��\/��k|�C����[�ٹ�5�R5]�b���>b%R�y�AE�H���ȴ��D���/>� |�h�-�\�az~����^�M�z|�^>/��៎Z��O�����P'�_4����j�C�RN��5C���恄�ݕ���Bң�^���ę�����e��aN���8���z�ǋ&:/�w�H�,�Դ�q�Wu����W�#ԣ��v���gz�B�?ػ�����az�՛Zw����c_����$��bX+p)�m��-��"\�V)��[�� 0>��"p�ݛ� ��N.F/��
ۋ2��_< �0ٔOh�;��+�㲅����P��b8<��kxTob,Ք���HxZ��2��bүG����.�V
Ho���wi���������˅����3������vtp}��x��A	[p|����o�Q>��j���D�-���-��}��,��h��I�=A:-0m�i�PR�f{
�z��ae�>��0�J,�� 1��#�orz4v���~pzÎ�=�� O~���-=���Ts��q�$�<yl��޽2H��6�LE�V4+�w�1n�BN£z�\�)��A�rV8���C�3��J��Y���u���HEC}�}A�59�(��'��ud���<��k�b��Y6#ޮ���R�h�-�5]w��""Ȱ}.u��3�Q�P��ǚ�=�T;�P{�IF�8R6Vs[��	�p�I���EF�6n Q;Od�f�N���=���߫� ��pwҟ�8�0�j����T�ѽ$=��p��e��9�k-�}�����0�noZ����i�\0dE�fֿ�}���f��f"��r�<��r�%��7��]���,,8����<��\�+�.kߥ�
�_A�&xHð�ᬿ��E� �׊�`��[��L�=�K�:��1�@Xv�*+�вC̉Yo��@+TG���l9 q�����1w"U�P2������P��M�(u�*`��`	��<aS��ڭ�\�=�Y�`�������/Z��N�{Pc�0Qj~k��բ8 ��򬘰(>Q�����Z����˾r�D:�Z��tn�Ђ�y�{��m�z@�R�����C�
�= m��	pA}_C�Kћ��o����S2�'F��.´����"+;�6"�o:{�0���ػ��$���#˼|�l]t޲�;��9M����ӂ<���8�"�z����z�(Y���c�����p�W�0}�f.c[¢��+�\��D|i�:���V�O|����]�0Ff?��H@�>�т�c����at�xb8��S?�F�]nK��;rzX,�&hS�Z���kIg�o�1U��Ų�4�)��� ��o�R�v�D6�>K��Z�'z��0'g�Q}:c����촄��6v�� !8�',^x�
����ЩOT�i�۸�l��d.�����n81�p�0�}��339�bu�]�����Ƅ���	�+��ɥ�N�c^� ���^;�[(F+i�j�씥���ؓx����V����;PHͶ��D���H�_O?�A��v��jJ�Ҩq����}1�&��M�I+V���1��3�i���y=�;&��ʉ��Vq�?��$�˲'��JI�&yv�P�SO�?��m��f���U�hj���˜FH�7e&���{��i��6ZP�4w����=;�%|W�__��ș�>Sd�i�lA9D:�۫2e��#��*��Rf������Եk��p�R؞Xgɼg��W��^�Y��s�Σ��;8�Gs��B6_��?�����"O۪�O�Ѳ��.#O����1������m�G��Y��~x�%'�� �~}8��M+'!.� @Iԓ!�Qqw�0+��AE�C�}���`H����g#.��`�-�&&Fܭػ����b�^H�8�p��˸�f�w���J�I�ei�t����W�f�H�8W��ލ��%$�KDW��f+�1��u�+ho�	AB�W�.��^9@��!ɫ��`��#�[�:��}���«<�z���M5X�Cp8͘*�5M�ZqA�4���+zq3�@��x�f�S9��i��:��,���\�4�m`��>�����aM��5�4qh���D�t�{���ks��'�������T�}g��h�T���H�{�0��Ω.�Z��~퀙{����7�EM7}]4/�jH��u\�LB3\iQ�3Sm�0�J!��Ձ)eQ�p��]=��h5۾�>A�w�E�����֍~b�!���%��%<�<�.e@ɵ���ή!YǉxÀE����ac�Q#8{Fm~b��BGa�x��L\�y����"��?�D��}L"�e3U�if8+wX�Nt�QN���w]9=4��ޛ}.����
�q��f�\|��|�B��#�{�h���J���J �U��MK�R�fHշ����Z�ܸ�zl���ֿ���C���K�F
�ޢY�r�q"n�H�?�U�w�ym�%�h��ZS*�L����~�:����-U�.���� k�)^V~�y���ӪD��7����],�|0�9�k�JC��,�[\�Mh�mv}F�a<�'X�����Jm	;\�v�����2+�6������½��+�3�� 3�� �b-%Ϣtu!��	���:�?�5���/i&9�!?͍Z��[,Ѭ &G�1�����w��R��*�6�?�"y�sف)z��[g ��;��J��wߔ��6Q�?��^o��w��}���41cpC-nj��B�C��dF�����>�(�D�� F'o��H����ΜFt76ͧ!���!�u�\��bA����^��h�Efu�}��f����y��{�DYb��m�>�֊/���+�k�#� ��~�B`*�yЈ�u�Z��A��m	��q��b�"��Q�q�9��&�^�����|�_�|�h����9�L)������h%���
$��,F}]�\l51���;���6=Z��e���a���4Sh�^,�n6�����(�fZ _���idrƸ�|`���E�T{�4�nQy׿K�]H���<����o{9F�˥;��%�_-}���+��ݒ�_O4�e��7V�u���
`5p��c򺝮M���~��Lv��6��R�'�"��W�O����w=��1_�
5��H�-��c��� ;v�=�t���ir��g�[�W��p�Rf>�J��L`�e�"����]�eI���dIY	�m�@۽G�ϟB����}���Ur�j�MR������!9x]�K���@�y
C��{�f�C�b��ʏ��Y쩒͉�t�u��#���dHeC�>��2 U���B]_)�qr=�*V��t\��f�%��%g���vr�ڗH7H�j!�.�_Q�E������jZ����V���(��*k���N$6�&��q�O�xm�(�s��6R~PU�L,�mWleF�u���U��a	7Y�+�Pv:eQ�{q�q�e�����8T˹=*�=tuey[�@p υ�Qql3�@@�z�Rh��+ܻ���Y��f�s
M�La��l��A�阠(b:35��tA(?�Y��{�����B���:묤����"dx��pU�p�i2�;B�`��ٙ���n�S��Ks����
�b,�>�n�]�%�ڰ��SG���b��$��_�'j�NF��>���${���j=-M���j}V���]����b,��_�c򀤢��~P޺�n��l�иEp{w��Hٌ��G�K=x��ݢ�۱�'"��-QXp{�T����қaojQ�=���E�_�_�df䋬@�j�$��Ա0d�������#�=X{o ��9r
 �3`��( Yg�bi�w)w���zQ��3�C�K��C;�Y��Ń�3c2w����쮻k)�n�V�nN
)H��O���fҴm���m�} �apM%/hn�1c�[ycR��� ������ F%�N�n�Al�m����]�s�2����i���:�P9�sl�z����~Uw�\���q�M���E��E��3����GK�t��s��Ӫ�UŞ�2�s�J%1��Zj+���&����>EKP��U�:���2��A�&Nk�N�(�߮��H,��_��'���)+ k1�6�׾�8���N��K(U�I� o�f��J�י�p���P�r/2пy�\���C���Fzp����Y�v��0Z ]�n�6eoq��C/-޶x�}�A>g�)��=���2����`�j�]}bق�C�,�����A�^o��EHC�v�8��K���5��x�D�wA���.�F���
y�P#�#��^�>6%�'�k<̗E�l��P7�UM��xm�i �F�u�c�#[<:�QΊx��C�t�h|�\
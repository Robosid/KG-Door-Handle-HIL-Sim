// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H=XL)Q/X%6UGGNM#\Z[K<P-H<D Z.H^%G.5S)""$DVJ4X,41G1-K%Q0  
H"@_RPQ;%7#T(%&.\=;/7"?'0)4;VWZK&:CLP(9G[[#;NM&"CS8;G,P  
HPY.C0#8IG#=+"%Q%]A!X9(_P<CH7UVRSGL5IG]G$&OBOZZH"6C#G)   
HES?^XFD*8LO!=LJI9I2@0;K?-J)SV2$):.+N(@!OE.QQ8,GSL-9;Z@  
H\7"_O\:)F9^]7YDS.S-?634X21:BF<:/@UU7\0T7*[QM!S)U_IL8NP  
`pragma protect encoding=(enctype="uuencode",bytes=3728        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@%CR/->W1F"*C^1ZA?M5JQ^G]-1![Y#.N\234WG[1)=L 
@RD*T^L<!T5 /^_5<-I+0/CY0!_,U@O<\)0#76KBUH84 
@QH6X W_(5P4R$^0Z,+9=XY"G2AN9HI])NHP66*9A*J0 
@0SRZRFPO-S.PT,8K%/F)S<HV)X79ZVI=;!BS(DJ"I0< 
@G1F;J98(K*+$(>#N5DV6/NX%HZ>F]4)1#+D9UMBFXAD 
@U?K'S28::1!U::EP)]Q-)0P$8J<1UXSX/!S6^8S<1LD 
@\&<=N*$5UEW-;4'BIJF&_)IFQ+TQI#*I@\7Y;>R_-44 
@(2 B4G9\GLMCCMMHS;;'A417$Z-'<6SVR7N1MJ5#YJX 
@U2'@?ZX6VTB$-H/@:[_\UU;OY/W;9S_9#8[:8N?$\X\ 
@1/I8KN<UA-.4\ 1X+-?;A*ZM\X\78"@WR%-/G:16J 0 
@JX35%4^QV)<7!2NXJ!-1CN=ORKG0@6[^U),Z?2@K,]8 
@*AZ:#&TDQK/Q:.IN%,9D].1B:VB)-8N&$LV\VJ1F7B, 
@/+/,\P/2P$EHTSK<P-S4L(XJ&$^D^A6S1U&/XY3AF@$ 
@?U6BF-V$/6C"]44XKU-YG EE5=D6,*7<I.*S"SU9X+  
@+Q^8J?4#;<HH;1\6B4Z-PACRW4!XWOS_N ./(,WL5T\ 
@W<KY]<5'_%)%=8Z%L@R.H[7E] F_GF,);+<6()?J-W$ 
@#%<\R-5?#*O+\VKF8?:]$SCO&@R&S'B"<$GK'HKB,L  
@C\]E!O>U2\B:(/^ @1Q2&3U+.D(R0HLEQ$\?./VX!M4 
@C_EO4J]LF53D%\XPWMHGS\OV!@<-NBVZZX]#KU;Z= D 
@8?[DT;71R82S9X3HT3_'\4+Y2)(*%F]G", W!KANXJ( 
@M\<O$#B-9'\G&.$*MO#^F0)1.A?8-X+ 59'@*2%%A:H 
@R5ZXSZJJ:X\MB]_M3\T:T?-NP\\W-/#_"&45]Z?>>Y< 
@$(34<2EGW&JZ_=E ;;LUN0W/0@!PF^<P2(C%?@=T;M  
@<5<0B(8  TJOKI[ $$_$<VO6,!=S'*WQ\?VN/3+G*9< 
@+N.>!-:U^%S97Q)Q,PKM0L6?4TED"G<>P%TBM7\8RFX 
@$=KV4KZ.5<'4SN]6]&LU<G\QS\E0\+A0IWUAB##&_KT 
@0G+"5[#,U[*<]W%>6V[(2%A2@.7:7GMMTOC<K;;<@3X 
@N%NCOP!:F!7Y76MU%=2WZ$VQ!W,QUI/,[QBJKM,,&6P 
@J+U+D+(\88/OVQ.9HH_2( 87IP(%H,LEG26C >XRF#8 
@\&>8>75MB9N"A.(Z[8ATEP[OBB+Q<7Y;TD2#H^<" IT 
@)!S_67-93-JVU6KU-#5X(+UGL9+1E&Y[+X0(6R1&\9P 
@0_?CO@D-<JM[ $RPE;X-?O)L#LP-])XD)5@/[54V>XT 
@' <GS_!Z3"YC_7NE?%+U2\<HC/0(%9]K33<C/089=H, 
@T0E%>*W-0_J$1:'>//]&:/__I:!O7$+4+2.@\"L0P/4 
@%=IUNK% +F[,#^)MZ<_$WCWG'7P[O\2(:FPKNGF9X9T 
@P/2B_EUX(U6J#?"LKD>;5 ;0L"?.5>6@=$I=/KO_]"$ 
@P0)XL$?Z#,AH#P9?!I76SL)<D[&1F,JVS\AWJ01>[CT 
@CZS1^=R0OR<DCF?G2E.T1<,I!5O*'8C6FAN_=7,-6=T 
@96/X\ST=U_86OTU#OM#6!-<^:Z[Z$9$K+KK:07N#R$H 
@]8:V6,; Y#]8)W$'HK"E3$L+^OJ#OZ;A*T8TM*D.'^P 
@Z(_T)C0&XF+$XF5E7SATJ4E>K@X=55XLV/#TB$7=H_( 
@ZW"C4'&V0;],^TU9*2,K7E?>.AH^+4A.;;["LL['F#T 
@J/%_KW1F+OZI9:\[5Z)B(K1G5MAMP*-?U&@N%YABVF< 
@8<ON4KI=VM[GBLRDP6C@V(D&I-;:=_S^R;\YFV$W('8 
@[WALG65RU<MBNL&KN*XEK6$SCJB@X^LPXKVO@0C[TI$ 
@40D3[_+NLN8I>:TY+MP8N.0I:7"-WNEF$M9!VPCKO3T 
@\O#23H^EKXZ9@?9;!>.\ S>5B<_$R^[F9FB\6C>2$U\ 
@.KJ+/CE.RM)5UEI*N8@#CGR+F.EK96L#3?EQO],'M T 
@/'L$=/8*PE"'7GQ^4YNSQ7!7&$$'  XOTTRF[Y,S!&H 
@#U4]VT_.V> S-;?P:?Z6)?@^2J_EVHA!J;T;H#: D4, 
@CN<6[D.2(GWH%8.W'F[X)%M$U6'X:RP:[_8=&U14/\, 
@BSIC/^?I2.4_YVCN]3-WEVJL;C9M/&C@>-A^P2-?'6< 
@E0HV=7D%U9WF<EES4?P%M1MJ,AV<F_"BN;$!$7_"#4T 
@.Z2ICJG?OU3SYF(FXZ^6MZ@NI(.OX2U"U>"$\,E 6.D 
@1H]'R<I%R*8]:84_"B5#4(2Z6ZM=<#01#FY5$6I+\(\ 
@5UO3%Q7Y2U.-AS7$A%]1!T2%QB<T'7,NF__,_ ")00L 
@<$2>IU^"D'OU\Y<J\MBU2W%?$S\TZ::BF&T?D\4_)F@ 
@DXHT:,J;'I*[^(5_YC8MJ(MJ9($1/A=R65W/")^=780 
@ 1L3;50SSEBM4QH.]B\B;=4>J\JH#\3_-(?I3PS@-VH 
@;_ID1.18B,A:JRV4!6=E9TY%3TBZ"01,US,#EN[;93P 
@*^@0>!DL\"!E -L8ZPTSR][@87HDA @V$ZXCE= >#Z4 
@[(A1G6:DB3M_BL7E_$</#J$"C>?%4ID3 F^.+KW$?OD 
@6?ND'AJHP'(N;K'W HJ%?OH"$(9W5+57#<C*K%W;UN\ 
@.+CA6N6(EG.\K%>Y(E961R17I<<H[TL*8SP5CAZ>2B0 
@2'C$#'W!LX#/IJJ>O6#BH_<AE8GUYB?#3Y#U0#E'[(4 
@<]- :BA<.1P R._.9"EGI_\RW !]1^L[^V,9(R+HH&D 
@$QYKWUE6O>E E27QNYVY_Y?,=>&\9:$HK.TA-XX+1A< 
@\J>P7'2P-;K#ZG7)PH0NIP2[P\?D>FK4CY%6^-3@7,X 
@XR^FVG^8_Z4 /VX#CG5M#:S7]+T.<)% 8 IN6D<H6V$ 
@YV H9-V7'<->B]S\"8=+W1',E@,>5=V*C)5'7J)<Y]8 
@$LU[+"_?76D+:B?)1ZN[CCFSZ91W_M*/._\L3<4;LO< 
@UBF/31^_Z<!B_L(Y-DT:3YT&\GPN'NM?3WOZI&*YW:$ 
@GG)3=ARSX27BS,DN%TJ-_!#8=\Y3#RIODE6L5#;AQ00 
@;G;?E%+4/^]Y>5C2GE"=?#1 -Y1PJGH4LS>@O$!=NL< 
@4H9,^KF;\@1K29[IZ1?F,47(>+@]V&!IM:/3N!PJW,X 
@(\GL)!A;V6/WV=<.(=;%)P/82^=<ROG7;W =2]T7J+P 
@E-)]3+^69[<T<_#S?P9Z9X1Y(>0J(CY8$0]?V%-D2U4 
@ZGF[E04:J K^X'I$)3D<XCNYF%7B\S[_'-703[![*NH 
@#ZAT7J/S(&/5,TGP,O#S#0>D7%CGM&V]X$*,5'RXW[( 
@?4F?<?*_B&CQ HXXC&6GFQ++W5$:/.4O=M^P/6=FSXP 
@VLU5@$E(,),,<](RH2-H A5D.RY5P*B\FD1+-MFQ?5< 
@VRS=4#Z$E?(H<"]R@O>-.E1C%:BTSD=] -W5O)NWOS  
@,"#^RD:DG0H6_/S*/" ETE*G1,,,3'TEF*U%#1^4I9H 
@M35BEIF% S^#JKI-+J>+;A*2IW:G;BD!KM]6.N("TYP 
@6#% :$UGPT;R.;!O?7H$:._#HCLR(<Z6GXGH5UE"NW, 
@$=GV&:;F]8>#\6*G4>@?%7/L-"JBJ<;!(LU:((:A[$( 
@4JO1XD^Y9V]97_I\F^K$4]_7G7;FE  VS<?%M7A%'Z$ 
@+TW)RABW<]B4H![B$$/.# AI_E4/[WIF['C$U8@?;YH 
@";!"X^%6*F.D0@@4VXR1GAFJ^%)8#(:3%TS"^N66ZGX 
@593H7OSR[BFL9)*344!A65*!#PP@#UZ+DM+<_3G,+8X 
@M[;U!.9B?Q+)&AN\JXRIC^54*]_6.>PDQ\;\VM(Q6N( 
@C1*75]Z*WG1&)'H=:@6%Y\,70=@/34>L\=B.L=HQ6)@ 
@\#1W2$Q$[)\>"9(+DX]1*@]W?M1\5^62:DB#4VO$Y]8 
@:(E7-:;(NZ;4R9-ZS3?'G0!B? -,^]:H9'/NS?PVG;8 
@RH7*RPG,;O$UZ_EG\'EN$3%[N94)S8.G 3&MX(;546\ 
@$1W>624 *!?Q#:'WG2(36<DE'!&!+_#O(?2-2MQN4'4 
@<GI" 2(@-4+-K(PK.K_.%Y;V,ZRE 9VS7#V(>,L^P?P 
@M<^,[KH5TGPD:S83XRWTO;!_O,^Z,Z&"H#,.U\:4<2$ 
@,6!?3C: G Q!0*N/?<*E453AKM_\6TIJMJ#652L)/.X 
@T^+R%N[00^+[58I_4&M;/^/6_;3N)V"887$-:PE(EXX 
@V?23.Q9&MBPH:+'+B>WO3R[W4V&L6"5F:R3RQ2U#1I< 
@^$)":<)64"=.EHVG14CU/ACE$'D:OYZ)Z@V?3YB+R5\ 
@95QBR]45&8[=;T8GIB9V%(W[N37..=>JQOV=_8+HG[0 
@HYX?D>R/B SXT_>I&#W>4*)0F4PW?6 .+*E+Z#[?:AD 
@@8E*TH=[)JKC\7I19NUE&8E(O;'5$4 G>\T=!@/67^H 
@J0)8?$"UR9P>5&2YX<R=2P^CJIWMYH@2SJ;/M'<KVZ\ 
@MK;!93.&)TV3=52P*(:B2]_2L/=>ZF@2/[FAN24$'1T 
@H^<C#U%4G\^AUR>)PEC*W/>R!'DJ_P&9V>^:Y<_2"%  
@J,9BTZ5?MV;()5JB"*^KCP $>7W?+,[LU@\^UK$LW>D 
@SK#9:)EI;&];]S%2=H*>W)/YP@:79:-]VK>1E4\)RD< 
@KK#$YA[(!J3516I^4V)7/G+VJ7-"FA&P@,],I7+G"=P 
@KDZ'"I]7;V=]5[&EB;)9Z,L:^9Z&-A.=@RN2$=1,E,8 
@!KF^\]RA9[4&CE'.BN,GCUGB!%QI,?1BMPF.FM*M?5X 
@-1[,ZO?_S]>(\9J-BL, I2%)U#'C/9BKA&HPNKXJC6, 
@L#C<K9P/H6_(%Q,K4U4%T%V:>BC!:,;74%R[YY,Q:^T 
@VBX2\U#O^GF)SJ'AOMM\OZ5.(O$#4"T*UWPC=F?1HZD 
0/DW]SD1_X*%W^=O5K*)[K   
`pragma protect end_protected

// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 12:34:41 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FNwwd91WUiszds75Fo2HIhMChUod9gUU7akwzp8zPyFxueZwJifnxLlKFB/cGyA5
F2xsB4jAmmrgWsAOA9K2k68lyHIZ7n7levNwSy5ZJFHOf0NbISAF6qrJkA2c8dhC
CmBcxweMDmZQHGJlmMmlPK19TA/rJYG3bH4/kwN/6Zw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6464)
9kzrhR95WeCSLderd+vSCguxUiHC+kC6u4nCRHrZluj6f2vTyPLOpxu3/tLKyjPd
XifSSSGC0wH4/0OItPi+4qo0qdBH+/pqRKM7dCRbgDhNBEBm5viuYp+bQ3lPnjOY
avDHF4CVdFjSXEUw258UF9onue/T1C9FTNaeSE3nlwiLI4I3KWQ111B6PbFoWa0E
wPjZRb/pR9jAIU7eqPMgSFVqBxnVosZSZN01SsOr273ItjIhLr0awiZYzLhF32LB
1zCQWdFaBTYdp2yJ3DSZVMBI1rOiTAc9oWSxcToDqr4DOJ3kO9QoNpmIbp63LNl8
8O5qpvmpPxAFmUd/SL3RP9nrd2gKdvuF5/OVsrihxfxtqI9fVrZsKRicIRFzylMl
pR3nhjEmTVE7Ymw108Vze/AUvnY8DoNzVzXTfy8MamlTxkQotfYAzlznL0ceDyMJ
lIKzkWo4DYOjF/VUuIW/fmJni9gC7Xjdojsa1HqJxAuqzZkUOZN8c5JpdBIVcB6A
UuQiwoDD7g4Zsm0irIdRFbttSwPAny0iONZmZ7Oim0nx9Y/DYKfw7+zq5ejZgtCr
JXtauggyatU8N7Ax3aaW2Bxkm7sQ6bLYtMiFSYtkILFSDsrR5495s4otTHt+12n7
y4rHuLDdlAHiuq9jkIHHXj7ih4UJpnxnKnf4Y248p2GRG7nxKUVmIRc61KM5SvAe
CFMue4CQGzd2sDKl/IhZk4TwdB3byExgAhEoFUMofP0Pymxysiz5Ke0DhCTD69TQ
pp2K0DzJxCbnICPrilB0AItay9dDEnsOFeIsrkQ/edO/zG69EO58E4b3GCQBqFQo
xgtWJCklGHiMSQ/bsLO/bSQ7xQMOGAq+w4bJ59XVCZYn82zmIz8+DL5zu9qshDGb
mjQibYRmwn77FDmQeb4MQXWmuKVm3XHwRE429mos3zLkg6HBVtQwff5W9YlQqKi3
FLzau+cF+aDbVE7h//bvxHei5NDQOTqqT0etZEqOE3vJKgnrZptymk1g77xBfdYK
5hiIG8SHd2yRYShb9VL2bgJmiQR9hgjtKTapyMCnoazkE66u9MB4IlX+VAaoebxj
SDcoq+rYNxY04bylT6du3iIRUIPgtEXImdhsSp8YMJ4AqLrCukNtLoTzFJ1abzgh
N85W2PoizFMG8hd8pLmd27/iAuYXgZJ5WTKWXJNGFilhna98FPacqq/KZ+sa2yVD
DT2eF85bAxyz6pTT1ykXVXsYGMRvdmgbTwvBaE5MGRoJc0kgSf1CS38gPRBT1v+9
F7Gu6t3OGy742bKWlVKYtCCOb45Wi/qhM0c7MsBUvnBY8rMN1uNfu5o621225ImD
N6xyUIOgJokdzBFi2YpiF1hJ4zIFuy4u3DMXP2p9z88ughDVyNzVEpwvVDRg//Qg
HbAf64428nFqvFdHArQdUhFETXVHKzIwnw6dn+r+lLhSLie/dTGxd9w7GKtZ9rS9
BvdyisNMDnwQEQvS4Aav+wEgb9H+DL5hswzTxKCtDZEtEW+VBp7uEtKtT9gm/zAh
rOrR31NjPdpMKvmmRhbjfunPAQQDFiDLDDg6CiysYh2nFFwaEW1705YML7+8O8HC
bKStbXkWexLAuIneXBBsmEwq8amt6nYGuj7PXRWGIQ9UERfG3NN/tIKG/xDHdvob
CzcpuNW6VKF/akbvpJFtaO27GgFCgJl80kCJYZF5bhqAOxXoOaWkehcfN6Rhkcqr
XSG42QzSysHEKdfA3ollazeWqC2tlKS/QA1p0+S3hnmaGB6ZiwGooPdKWqgEDkT8
oBAWk4IotsSu5fGnNOSatt8OkSs74xU5vWmb2U8tkE6EiuCkJOn2ZCjE/KUmToIm
gyLQZf6RFknQ2tJdoZSbfuzwkbluRsSikuAZLxGqnvsI48RlFOwDziR6C4xrtGoH
n6/Lhwk+QDVZl4ee8P9YlAC9QIiB8uIkiVFphgBHjz39WvUPPghT2F1UpUPRiX3V
HVMrTnxiZbEXQCq/onWdz1pfFVLyHN/TNQpWYWjKtgHgi4X+YDqwaP10oI7ixBd8
B7mGcoNCyj9nGsLPx+bvPTIu3c41Gvda41o5uC1z9su/4qTNLn5U13V4llLWQxnT
qWHhtRqAFmM3YkSv3g3rtIV0jEVsVplwuPTqzKLaH3S7IPr/7qDzX/zROW1vUSC3
GX7JvqFQR17NAU9M0V04ObRRmlKUStuSW2yipMaLqu4SHEKnofIFxdUN1bno784p
bZUSP8iTG8HV+RjSzszJclBfumj2DSZy3RGA5IRbhD+Q5DQg54QYIoGAN7n6fUAJ
k2zUnSLalzG1ejVBjp13EAviRLTPZHWDXffv8ebNIuIGWTfR8TpgS3UtM9yFjF4y
5nCw/RJXpmAyiRpr4iGTMOVMTxAWXDm5DeRFRkG/TtgAGxJ96HzMMsvckiH7gDlX
HZbyt4lJlDCTB/+nffCR2oI9T0pAjnoDFMaxgm6D7j18olnvidL2s/TwLMumLUuA
dTOs4AMDqDfUR6Bwl32ouwXvXdIlNPpIpATa7ZMCN17ZiXhIPwEGYEdRFxVA4pjO
QzCRiE7siAtCAYFbpxeLn3+DPcUsmIkm2FViIaDR/jSmRPQupS2ZMeEDtadNgTXe
eT6tsXeb0/D3ozrqWesxy1LZ4QCYepH/NSN2ggVjpnaNr5TeQ0I+JjG9wc33D7vJ
7gvZWEXBctPNtrS0/b/cbxlyEVMdyQTwUjhTmoEQxeJcjhkdwNn6ry0CwpS8qwB6
0qHHsgbotupO/cloKdlyFC9HpQHRe6Rn7VGfghjF5OJP243MfelzORMvufGk1Uor
X9/pICnfHIwfMTdHB/Hl6gNg/s/6mK8RAUDAkZ0Luk6w1h4FDzVMKyjxytrdZodA
hNzpis04khBQzOVdUewP+muKklgotPDW4bHGdgCHgj3AMGc7exh2rKTnns9UoEsN
4dOvLNqJh0ImoFebtICm4PBgCRBdltbyvvR0xKWUirvyibiVDvl+U1KDnXa2kvvY
rwYipsR2e5TV6cLTF74plJUDmMUIPt+cvM8KffQMneuERntFNfQJ8IUz4oGzAC+O
TQ7D2pQOOZcwcX05vcArTfDfmXuE4y8pxGymfgftt4E1LLoGK8ZB5n5VgUA3Ux5c
VVxegd8qu0AFgeu7CkarL6zt6b2C0HbvxwvGL6Kxn9BvPlSjTWCzL8SzImGBYN4R
CL6g1KLMel1nnKLdRMbjI4Zyg1lAoW1uqHSLbG+rS8uK47YHJpDJeZfb279BCNzg
QiNU41Qno9KbIkDCxEylFpy06LYz3fb78McgddlanrNTigr2uuE8LnK50JZcdu2k
2dZtCDlilmYg26kc8+gYPDFlyZe1g0oRSckvcEzoJvPFxPoySjJ72PPonL+vgHXW
bGJPLc7vFX9dNypFK5Oz/CjCQGXb0/dKSinGp/H+4rKx/wRRsZS9M3OjeIZ6B0ba
y9Zmg4VV1pYaSU4jCJrfpfYO9oNt6e53Rc3rrl/Z748cfXJcasasD52NEuttZTDx
0e1BpeuYHrBCnykpNrTdZoTi2R0aSY2z/dEkwocjjCz3JJPZUPVntBGGis9r5tu7
OhDGD24iMeTpA0xSE05aXxBJdqX9LVrJjFprnNA3cQFc4FdH0+rjNsbj5yEuO5p2
Zz4ftLQ1eoLqwEXK6F3oHVYBEjDHgAk5f4qY1x7sKzj8+tfe1XvT4sRpoCec3v2W
w2lWGxGOMWqRSMgz4zkR/QT5oPb8C1ZlL3TnM4WsTWKfQMa21n+OHvP6QCMtQQGD
eyBI2Z7Lj30MbJ0m2LlmGUMGCZSrb3jw/o6g5agBWpk+ANUmn13FkGRYW/0Z/Lsc
MEICjXQ4jjIaGgkjoKMfOAv2ppBi6EQIK6wf/XhpmVnyyUMHZ4/qYDKiPWsT/xwr
2razqGRh6QqcS8y6M+NGAeAs7X7foAvWa1xNj97t4YKPQan8iIxOkqAl+EmDvFIp
gSRQQMJc0wB3vr27gPI1PJ3ogSQOYYaBY2fX3NhDXCpWw2yCIHmFpLOBPRjFGXYC
WjTgdrGu8CuLubyCyKbLtjs+Y1fGYpiNlK9oZT7HxuXM7gtxmXtd9m5P/DtcpOmk
olL25cE828vyATCkr4b5o6KDa7dz66ogyO4fqQJ8SuE0FTVOLpAN8BMFiGYNKjgI
N8NEp4kLcJTZTOPmezAm46Kyt6K1YdkmYqXzKO0NuIebuk2/s0O0obk+9R73UHPJ
cSyobanqf2nS6jgBDYmh4CZh842Xtk2qJUCpEvWkznLiqs8qO7QhLdEMP2UPlEoO
r90lmzm4WJTHUrsahqRhthcxrruOCz+brozA1OR3ozQ7OKjJojFzyOBkNdIhXJ9J
7J2v/Lk7OX2Ky2ltrxVz7NLHLF2EPYMYO3pZJAVdlpuw0SLrORKduoz3/O4qZiRR
AZRkPPVeuXdanHGhTGZUbCUbpjKsUzsekhnBzruszFJORp85HZ9FgSFfASmBNZSy
asgxoDrkDa4qXQ4m1qutZi6lIP0eA5eQ2E7Tx94Z2ht4Z4HPmW+4+VgVplIUad8i
q42B+taU+GhYzLIx0g3c1XHMG12Tf0QVE2XAQndpZ4iytDmzPK3/BJ39qfafgdUq
YM6KUyYOZHBQhPp/wSh9+Nqs8NCpCqxXO/IUebjEZYg1mHXWH+IAGmupkNIwb6G9
AYgCVMX3oquRYFr/jKV+77kxo5bd+9G/FGUsqSp1ypgyr1pWYA+tDkHizD4Kj9bY
4H/4mEPUbQ3/LzbP9MF+cDlgo2vOVmaX0Id1cqzgp7syCu1umrQeT4JFyjJyoaxA
7/5MgfbNFIbMmm18HzC2E1oc2ANQrw8z/KC5QPn3vVdy2F5i7hn372uvHGRAAN5a
1NQ74RiG/z5mOPTGhBE7n5M29Cu9qvRON9WRaC9SZ5EFA/7xAFKKp2pCXwWyUY++
g/FYXZZhx6xwFFAO1zESw7zkLpMrME+CM1DiKJxQLEj1aWPyUbL6poAeQCLU8y36
X4mrLmaBLgGXcXy/70hhc7e79WDNFdld90boj7K7cLF8IufyeG7TJIN9bF34CmK6
QH4jr6C7u0CZdWta5oDYS36cXM/TMPicPcRe/SCNZ/ImkE2nLqhSdiX+zxelXK2y
cSuYv2Ju6ZvtyvezJxQizUf7THBOmOI03O00Lm4rCkRuTnjak6r+URTGLjTBSNef
h7fac/IG9yDrPx2bIiQeMn9SFS6nBQRlGm27MCTRKioR3ipXSAq6VuGUaM4ZRl0t
gIUZvQGRIvz3HuF1N0aPM+28wBVL75uuXc4BjpG8cbWEB3xFcCMP3K7tqdY4jFD7
+MtqyjYtohYMP5tS06XqUSC4kIxk72RT7gSbAhxdanHXPrfG3VAvoYNEHPniylmd
dZBf7J22vtKTr8nWZKIXxFtMB5gVFizkQxO8melS7zUWX8S09pYGjHJWkVDq+wcP
EmeeVMiWnNpFHbIlpxEWq2MGp1Q/+y0c30INVXkBLc83TWlkIFIilpPk0qIsMyXf
6A/tC5S4wN2qwoaA/k01mmW9jYeHSG45TU/eWxo2kOS6IGF65HalYb7/IXXAi//C
khLVyLJgpHF52foqhJvMV/UAnRcUItFXO8ysXXgkaQ9yfnGMbEH12sYmhJpEE/rd
Z9GbhkxpcA7P4RwWn8ARFx9IxXBnR8GfRBlsH8XlM8Dzg4OnleuVp4ePM6JUe3s9
dT8yyhQCn6mQtL5Pm0mnM9gwle5ONcJh1+qfhppEcKzxGoYa3EjzJZDpHrc7EyiG
DPYaB+HeCU9ROnP8ApCUaEQ/rP1f+YisqNUr45L8vRljpTIdCTezRklN5ZX70UTH
ygIYko5W1fvqPWJh5ufHyPsspt5pEqcYhRgEnrFNDZi8AJJj2L71MZ+MK4zQppEs
O/EjKKaIxpCQHv5a0SQ41M1rghwNVryvlFT7hEA0qlmw/ViBSiGHHstFYVyRei0A
PWuRl5DsqZFpgBtjH5Wac9cYslHoJoaH1BHAPUpsmufCgQSdQQfoYMmrQ9jygRIj
HuqnzkBTGuYsuiy4lp0QeBfN/x1Wk5DcJYbFCT4zu89EV3GKLOcfU62Rl5UK9obO
CkAuLLNgDdHmZAk84XxNVrojAcqqZWdtGYJ2Q8OJCbhpe+r3G2L/dHBYnxthDjAP
deheRwPS8B/EuNGWzYag3yuNqIyQmfaS6EJQn5puEGUgcEiI/Q47dM+0WEf1/ct4
FqoSYHKiTtxkXLQ7S+ND1AnnTQrjVyLXn4YchzZkJQUYzuUGHeYMyWfL0XGbPzAq
7GK2IxDp9QdWO1HlNRKHfFLaBX40mDvCtH5vNwZ67fuxGNVY8at7suj8fVEe+MvL
68gXIKByIRh0QWsYBOLN/r8Xvc4P4uvblPF3Mqht/5cLeC5JjEev3pvDfQAvP1nM
Og6j9hhS3bk3gxYzV0jEeEK9uZurqCgeL1KoYCAIcXIKD2CYY1b+ku3f2Fssdlsg
kCJmJXTy91k9BB3d8DZAf7eieH395mwxebijTIexmcYuhFIsr9Qai87exCD66a2b
eq8YNDLa9I1/BTzSFDvA+TaMXLIGIBQHiC2E6HvJg65hRaZ28w7kk8lY9WZYFjm6
8fi+aV6EOV7z0bMCcM5+ZTswzurand49+HB4Il11DtbNvK0Ia7vcTgwXYoweUNmL
vap/m64GQJOyNUoAVFE18SakcfNiBszb9VXNfjpyl/6aw8b+MCtX2Cp4Tv+eKrbI
T/abCzPxDDz1EZn9Z9rBfGC5dpQbn0f6n6IBv/pr/i6fCGk0aH7e4QlE7tPxmucL
ZB+PbG+DBTsRB2thQBVXAm2IJ553haZOzJkbF4TWcmMztsAlo7QduWWCvg7aE83o
YTld+sHe5p+0GJv5f9GVvtcvWb+tzf9jg3VHRjrUHht6yiLk2uOeGUcdjwKlmEPz
y1BgyBoekZaPEwzy6KZiKfe+KrypI+bY29EclB0xh4DK1xN42PGPljHpQWxW5oJA
pfvcwCSBWDFLZB2kfcSoGK/pqDT4HzM/b02BfXzsdXyEYO2wIxXASIbO5J+0fqn3
fnwCVk/I/seK4z1SjRMjzsywPSqQaIuPOfLR5bi+blATt1VsBf+MCWABRAEAtM7H
dKeOY70/TxAbdz4/29/fNCXk8pUxqCAOpY4UthDUrr7lBT/tMX7TVgrkZxVb7V0v
UObnzuxcJm4jl+RCYQ+P0oEd6Ieh3R5qN5nZ/UY3+e9PQOJHSddSsJFndTGOyLdx
Gx2MRr44xd5HjHG/D9g3fSbupCQRZILi+4p61XHfyB2iryGZCuUQiCV68jPCtgJ1
F5MwVFdxquYq3XYQkcr4ifoT+mtzThWq74PePuku8Yi0Cfwa7uHEQf6Dd/RJPEDs
MlPJGMnv/uWndEuhhBTZuDV/2lkHAH7Xcg52funuLV8KDKZ0Ri9IupUSfosiCo/g
2XeJNatM7iXCJSkyMu2qVwP6qHofGCiCJmlzU9G6yMBlzrimjCZqluxSVIsa5tMP
x7wLAk92NQug1ceBz9uNK/BygPxg669Xr0tLBQ616AmrAVAZvfH5NlLPytezvjmW
aV6VFhuEyMqRxLt5g86GiSgCrZOoutlc+glbgpDU5NxIyZdlJOjxEJCx/qcxCTUZ
NkjrEJUPQP1CZPJc3CAzhAH08M9du67fUs00z1+TTmn4XORVZSDLmb5Tor0yg77P
Px9WS+X2q+4MPliACrZXE0G9JcXFNDyLbHB7Pqyws/++Z0aiV+GeWuf147N7981j
+VNTKNNf0nne4TYVZ30iBZEoTjRzryBJzZAHAidi8R9VsMh6z9zrABUVfjXmmT9m
lxRO/2+oWY7eVexXQcHDgxDi/kv/rcNroOac4mtmTyeaO2A99oN4hjoDxghfrCYF
vDgzcTiO/iVN3RoWZVx5JGZOUqeQJcR1vECjRPKvDtvaP1/gdVDU6D16Fn3l+9qE
05miiom1wJXNHNSA3FcQEOeDF/kksC7/xhfpwrtJu+y9OqM8niZFyT7l6Q78iiPR
topq+l1UqjDn9gt2JOBtqwlbSDHmArcJYwb6+kIH3fYlm9BRH3hDrDQbzOFCym8k
ZBuGi/KHD10KX4ptPIrZZRe6h0AMbcLVtUlwvJvaGvdP+5cYY0AxQxpcfrsClicB
RE7aUAXQzjA3x2VPgIdfqGtYFUxJG0X08vrx90w7uVR9feYVIrLZnlkyYimLW7UR
rhdtFAMBnLkKUvfxVktalhd84KB6Uc8oTgPc82kMqRVrSB3gsBT1riT1SJIK/OAy
NrQ0Z1EeKRzddTFDQshI7yxhzi8DmRnzjeasjJCGId1Jem8YKXTZeUJPjWPgtw+r
nVMUq5DErdsOv11Oi+7qp4asteffQAz8NxxwJu8Dd5k9TkddEoXHcu3ZBJ3e+j0q
wIQiPksckn4ekHji+OdLvpeXfPxjjmMGZ4T8wvRqXsYBwidXdRDLiFisLm/nT1WL
ZG2wVG965/DxZMey2G36iX/RVo/J6vtn7rVwAwOHVv15tE1A6LMhzRwoy0w/2QyX
5xsVq4zpWVDcE1d9i33Fjb3PWInDtIeiccwnNeetmaZLt15hgKNWwMMT+/E/mjK1
Qloheuvt6uoXn1Y2cdl7ylxYwJ0jt/K2VZg3sPmiyc8=
`pragma protect end_protected

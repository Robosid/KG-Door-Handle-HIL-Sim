/*Copyright [2018] [Siddhant Mahapatra]

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    https://github.com/Robosid/Drone-Intelligence/blob/master/License.rtf
    https://github.com/Robosid/Drone-Intelligence/blob/master/License.pdf

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/






// qsys_top.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module qsys_top (
		input  wire        clk_clk,                                                   //                                                 clk.clk
		input  wire        reset_reset_n,                                             //                                               reset.reset_n
		output wire        triple_speed_ethernet_0_mac_mdio_connection_mdc,           //         triple_speed_ethernet_0_mac_mdio_connection.mdc
		input  wire        triple_speed_ethernet_0_mac_mdio_connection_mdio_in,       //                                                    .mdio_in
		output wire        triple_speed_ethernet_0_mac_mdio_connection_mdio_out,      //                                                    .mdio_out
		output wire        triple_speed_ethernet_0_mac_mdio_connection_mdio_oen,      //                                                    .mdio_oen
		input  wire        triple_speed_ethernet_0_mac_misc_connection_xon_gen,       //         triple_speed_ethernet_0_mac_misc_connection.xon_gen
		input  wire        triple_speed_ethernet_0_mac_misc_connection_xoff_gen,      //                                                    .xoff_gen
		input  wire        triple_speed_ethernet_0_mac_misc_connection_ff_tx_crc_fwd, //                                                    .ff_tx_crc_fwd
		output wire        triple_speed_ethernet_0_mac_misc_connection_ff_tx_septy,   //                                                    .ff_tx_septy
		output wire        triple_speed_ethernet_0_mac_misc_connection_tx_ff_uflow,   //                                                    .tx_ff_uflow
		output wire        triple_speed_ethernet_0_mac_misc_connection_ff_tx_a_full,  //                                                    .ff_tx_a_full
		output wire        triple_speed_ethernet_0_mac_misc_connection_ff_tx_a_empty, //                                                    .ff_tx_a_empty
		output wire [17:0] triple_speed_ethernet_0_mac_misc_connection_rx_err_stat,   //                                                    .rx_err_stat
		output wire [3:0]  triple_speed_ethernet_0_mac_misc_connection_rx_frm_type,   //                                                    .rx_frm_type
		output wire        triple_speed_ethernet_0_mac_misc_connection_ff_rx_dsav,    //                                                    .ff_rx_dsav
		output wire        triple_speed_ethernet_0_mac_misc_connection_ff_rx_a_full,  //                                                    .ff_rx_a_full
		output wire        triple_speed_ethernet_0_mac_misc_connection_ff_rx_a_empty, //                                                    .ff_rx_a_empty
		input  wire [3:0]  triple_speed_ethernet_0_mac_rgmii_connection_rgmii_in,     //        triple_speed_ethernet_0_mac_rgmii_connection.rgmii_in
		output wire [3:0]  triple_speed_ethernet_0_mac_rgmii_connection_rgmii_out,    //                                                    .rgmii_out
		input  wire        triple_speed_ethernet_0_mac_rgmii_connection_rx_control,   //                                                    .rx_control
		output wire        triple_speed_ethernet_0_mac_rgmii_connection_tx_control,   //                                                    .tx_control
		input  wire        triple_speed_ethernet_0_mac_status_connection_set_10,      //       triple_speed_ethernet_0_mac_status_connection.set_10
		input  wire        triple_speed_ethernet_0_mac_status_connection_set_1000,    //                                                    .set_1000
		output wire        triple_speed_ethernet_0_mac_status_connection_eth_mode,    //                                                    .eth_mode
		output wire        triple_speed_ethernet_0_mac_status_connection_ena_10,      //                                                    .ena_10
		input  wire        triple_speed_ethernet_0_pcs_mac_rx_clock_connection_clk,   // triple_speed_ethernet_0_pcs_mac_rx_clock_connection.clk
		input  wire        triple_speed_ethernet_0_pcs_mac_tx_clock_connection_clk    // triple_speed_ethernet_0_pcs_mac_tx_clock_connection.clk
	);

	wire         eth_gen_0_avalon_streaming_source_valid;                            // eth_gen_0:tx_wren -> st_mux_2_to_1_0:asi_sink1_valid
	wire  [31:0] eth_gen_0_avalon_streaming_source_data;                             // eth_gen_0:tx_data -> st_mux_2_to_1_0:asi_sink1_data
	wire         eth_gen_0_avalon_streaming_source_ready;                            // st_mux_2_to_1_0:asi_sink1_ready -> eth_gen_0:tx_rdy
	wire         eth_gen_0_avalon_streaming_source_startofpacket;                    // eth_gen_0:tx_sop -> st_mux_2_to_1_0:asi_sink1_startofpacket
	wire         eth_gen_0_avalon_streaming_source_endofpacket;                      // eth_gen_0:tx_eop -> st_mux_2_to_1_0:asi_sink1_endofpacket
	wire         eth_gen_0_avalon_streaming_source_error;                            // eth_gen_0:tx_err -> st_mux_2_to_1_0:asi_sink1_error
	wire   [1:0] eth_gen_0_avalon_streaming_source_empty;                            // eth_gen_0:tx_mod -> st_mux_2_to_1_0:asi_sink1_empty
	wire         error_adapter2_0_out_valid;                                         // error_adapter2_0:aso_out_valid -> st_mux_2_to_1_0:asi_sink0_valid
	wire  [31:0] error_adapter2_0_out_data;                                          // error_adapter2_0:aso_out_data -> st_mux_2_to_1_0:asi_sink0_data
	wire         error_adapter2_0_out_ready;                                         // st_mux_2_to_1_0:asi_sink0_ready -> error_adapter2_0:aso_out_ready
	wire         error_adapter2_0_out_startofpacket;                                 // error_adapter2_0:aso_out_startofpacket -> st_mux_2_to_1_0:asi_sink0_startofpacket
	wire   [0:0] error_adapter2_0_out_error;                                         // error_adapter2_0:aso_out_error -> st_mux_2_to_1_0:asi_sink0_error
	wire         error_adapter2_0_out_endofpacket;                                   // error_adapter2_0:aso_out_endofpacket -> st_mux_2_to_1_0:asi_sink0_endofpacket
	wire   [1:0] error_adapter2_0_out_empty;                                         // error_adapter2_0:aso_out_empty -> st_mux_2_to_1_0:asi_sink0_empty
	wire         st_mux_2_to_1_0_source_valid;                                       // st_mux_2_to_1_0:aso_source_valid -> triple_speed_ethernet_0:ff_tx_wren
	wire  [31:0] st_mux_2_to_1_0_source_data;                                        // st_mux_2_to_1_0:aso_source_data -> triple_speed_ethernet_0:ff_tx_data
	wire         st_mux_2_to_1_0_source_ready;                                       // triple_speed_ethernet_0:ff_tx_rdy -> st_mux_2_to_1_0:aso_source_ready
	wire         st_mux_2_to_1_0_source_startofpacket;                               // st_mux_2_to_1_0:aso_source_startofpacket -> triple_speed_ethernet_0:ff_tx_sop
	wire         st_mux_2_to_1_0_source_error;                                       // st_mux_2_to_1_0:aso_source_error -> triple_speed_ethernet_0:ff_tx_err
	wire         st_mux_2_to_1_0_source_endofpacket;                                 // st_mux_2_to_1_0:aso_source_endofpacket -> triple_speed_ethernet_0:ff_tx_eop
	wire   [1:0] st_mux_2_to_1_0_source_empty;                                       // st_mux_2_to_1_0:aso_source_empty -> triple_speed_ethernet_0:ff_tx_mod
	wire         aso_splitter_0_source0_valid;                                       // aso_splitter_0:aso_source0_valid -> error_adapter2_0:asi_in_valid
	wire  [31:0] aso_splitter_0_source0_data;                                        // aso_splitter_0:aso_source0_data -> error_adapter2_0:asi_in_data
	wire         aso_splitter_0_source0_ready;                                       // error_adapter2_0:asi_in_ready -> aso_splitter_0:aso_source0_ready
	wire         aso_splitter_0_source0_startofpacket;                               // aso_splitter_0:aso_source0_startofpacket -> error_adapter2_0:asi_in_startofpacket
	wire   [5:0] aso_splitter_0_source0_error;                                       // aso_splitter_0:aso_source0_error -> error_adapter2_0:asi_in_error
	wire         aso_splitter_0_source0_endofpacket;                                 // aso_splitter_0:aso_source0_endofpacket -> error_adapter2_0:asi_in_endofpacket
	wire   [1:0] aso_splitter_0_source0_empty;                                       // aso_splitter_0:aso_source0_empty -> error_adapter2_0:asi_in_empty
	wire         aso_splitter_0_source1_valid;                                       // aso_splitter_0:aso_source1_valid -> eth_mon_0:rx_dval
	wire  [31:0] aso_splitter_0_source1_data;                                        // aso_splitter_0:aso_source1_data -> eth_mon_0:rx_data
	wire         aso_splitter_0_source1_ready;                                       // eth_mon_0:rx_rdy -> aso_splitter_0:aso_source1_ready
	wire         aso_splitter_0_source1_startofpacket;                               // aso_splitter_0:aso_source1_startofpacket -> eth_mon_0:rx_sop
	wire   [5:0] aso_splitter_0_source1_error;                                       // aso_splitter_0:aso_source1_error -> eth_mon_0:rx_err
	wire         aso_splitter_0_source1_endofpacket;                                 // aso_splitter_0:aso_source1_endofpacket -> eth_mon_0:rx_eop
	wire   [1:0] aso_splitter_0_source1_empty;                                       // aso_splitter_0:aso_source1_empty -> eth_mon_0:rx_mod
	wire  [31:0] master_0_master_readdata;                                           // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                        // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                            // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                               // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                         // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                                      // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                              // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                          // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] mm_interconnect_0_eth_mon_0_avalon_slave_readdata;                  // eth_mon_0:readdata -> mm_interconnect_0:eth_mon_0_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_eth_mon_0_avalon_slave_address;                   // mm_interconnect_0:eth_mon_0_avalon_slave_address -> eth_mon_0:address
	wire         mm_interconnect_0_eth_mon_0_avalon_slave_read;                      // mm_interconnect_0:eth_mon_0_avalon_slave_read -> eth_mon_0:read
	wire         mm_interconnect_0_eth_mon_0_avalon_slave_write;                     // mm_interconnect_0:eth_mon_0_avalon_slave_write -> eth_mon_0:write
	wire  [31:0] mm_interconnect_0_eth_mon_0_avalon_slave_writedata;                 // mm_interconnect_0:eth_mon_0_avalon_slave_writedata -> eth_mon_0:writedata
	wire  [31:0] mm_interconnect_0_eth_gen_0_avalon_slave_readdata;                  // eth_gen_0:readdata -> mm_interconnect_0:eth_gen_0_avalon_slave_readdata
	wire   [3:0] mm_interconnect_0_eth_gen_0_avalon_slave_address;                   // mm_interconnect_0:eth_gen_0_avalon_slave_address -> eth_gen_0:address
	wire         mm_interconnect_0_eth_gen_0_avalon_slave_read;                      // mm_interconnect_0:eth_gen_0_avalon_slave_read -> eth_gen_0:read
	wire         mm_interconnect_0_eth_gen_0_avalon_slave_write;                     // mm_interconnect_0:eth_gen_0_avalon_slave_write -> eth_gen_0:write
	wire  [31:0] mm_interconnect_0_eth_gen_0_avalon_slave_writedata;                 // mm_interconnect_0:eth_gen_0_avalon_slave_writedata -> eth_gen_0:writedata
	wire  [31:0] mm_interconnect_0_triple_speed_ethernet_0_control_port_readdata;    // triple_speed_ethernet_0:reg_data_out -> mm_interconnect_0:triple_speed_ethernet_0_control_port_readdata
	wire         mm_interconnect_0_triple_speed_ethernet_0_control_port_waitrequest; // triple_speed_ethernet_0:reg_busy -> mm_interconnect_0:triple_speed_ethernet_0_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_triple_speed_ethernet_0_control_port_address;     // mm_interconnect_0:triple_speed_ethernet_0_control_port_address -> triple_speed_ethernet_0:reg_addr
	wire         mm_interconnect_0_triple_speed_ethernet_0_control_port_read;        // mm_interconnect_0:triple_speed_ethernet_0_control_port_read -> triple_speed_ethernet_0:reg_rd
	wire         mm_interconnect_0_triple_speed_ethernet_0_control_port_write;       // mm_interconnect_0:triple_speed_ethernet_0_control_port_write -> triple_speed_ethernet_0:reg_wr
	wire  [31:0] mm_interconnect_0_triple_speed_ethernet_0_control_port_writedata;   // mm_interconnect_0:triple_speed_ethernet_0_control_port_writedata -> triple_speed_ethernet_0:reg_data_in
	wire  [31:0] mm_interconnect_0_st_mux_2_to_1_0_control_port_readdata;            // st_mux_2_to_1_0:avs_control_port_readdata -> mm_interconnect_0:st_mux_2_to_1_0_control_port_readdata
	wire         mm_interconnect_0_st_mux_2_to_1_0_control_port_waitrequest;         // st_mux_2_to_1_0:avs_control_port_waitrequest -> mm_interconnect_0:st_mux_2_to_1_0_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_st_mux_2_to_1_0_control_port_address;             // mm_interconnect_0:st_mux_2_to_1_0_control_port_address -> st_mux_2_to_1_0:avs_control_port_address
	wire         mm_interconnect_0_st_mux_2_to_1_0_control_port_read;                // mm_interconnect_0:st_mux_2_to_1_0_control_port_read -> st_mux_2_to_1_0:avs_control_port_read
	wire         mm_interconnect_0_st_mux_2_to_1_0_control_port_write;               // mm_interconnect_0:st_mux_2_to_1_0_control_port_write -> st_mux_2_to_1_0:avs_control_port_write
	wire  [31:0] mm_interconnect_0_st_mux_2_to_1_0_control_port_writedata;           // mm_interconnect_0:st_mux_2_to_1_0_control_port_writedata -> st_mux_2_to_1_0:avs_control_port_writedata
	wire         triple_speed_ethernet_0_receive_valid;                              // triple_speed_ethernet_0:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] triple_speed_ethernet_0_receive_data;                               // triple_speed_ethernet_0:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         triple_speed_ethernet_0_receive_ready;                              // avalon_st_adapter:in_0_ready -> triple_speed_ethernet_0:ff_rx_rdy
	wire         triple_speed_ethernet_0_receive_startofpacket;                      // triple_speed_ethernet_0:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         triple_speed_ethernet_0_receive_endofpacket;                        // triple_speed_ethernet_0:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] triple_speed_ethernet_0_receive_error;                              // triple_speed_ethernet_0:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] triple_speed_ethernet_0_receive_empty;                              // triple_speed_ethernet_0:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                                      // avalon_st_adapter:out_0_valid -> aso_splitter_0:asi_sink_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                       // avalon_st_adapter:out_0_data -> aso_splitter_0:asi_sink_data
	wire         avalon_st_adapter_out_0_ready;                                      // aso_splitter_0:asi_sink_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                              // avalon_st_adapter:out_0_startofpacket -> aso_splitter_0:asi_sink_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                // avalon_st_adapter:out_0_endofpacket -> aso_splitter_0:asi_sink_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                                      // avalon_st_adapter:out_0_error -> aso_splitter_0:asi_sink_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                                      // avalon_st_adapter:out_0_empty -> aso_splitter_0:asi_sink_empty
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [aso_splitter_0:reset, avalon_st_adapter:in_rst_0_reset, error_adapter2_0:reset_n, eth_gen_0:reset, eth_mon_0:reset, mm_interconnect_0:eth_mon_0_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, st_mux_2_to_1_0:reset, triple_speed_ethernet_0:reset]

	aso_splitter aso_splitter_0 (
		.clk                       (clk_clk),                               //       clock_st.clk
		.reset                     (rst_controller_reset_out_reset),        // clock_st_reset.reset
		.asi_sink_data             (avalon_st_adapter_out_0_data),          //           sink.data
		.asi_sink_ready            (avalon_st_adapter_out_0_ready),         //               .ready
		.asi_sink_valid            (avalon_st_adapter_out_0_valid),         //               .valid
		.asi_sink_error            (avalon_st_adapter_out_0_error),         //               .error
		.asi_sink_startofpacket    (avalon_st_adapter_out_0_startofpacket), //               .startofpacket
		.asi_sink_endofpacket      (avalon_st_adapter_out_0_endofpacket),   //               .endofpacket
		.asi_sink_empty            (avalon_st_adapter_out_0_empty),         //               .empty
		.aso_source0_data          (aso_splitter_0_source0_data),           //        source0.data
		.aso_source0_ready         (aso_splitter_0_source0_ready),          //               .ready
		.aso_source0_valid         (aso_splitter_0_source0_valid),          //               .valid
		.aso_source0_error         (aso_splitter_0_source0_error),          //               .error
		.aso_source0_startofpacket (aso_splitter_0_source0_startofpacket),  //               .startofpacket
		.aso_source0_endofpacket   (aso_splitter_0_source0_endofpacket),    //               .endofpacket
		.aso_source0_empty         (aso_splitter_0_source0_empty),          //               .empty
		.aso_source1_data          (aso_splitter_0_source1_data),           //        source1.data
		.aso_source1_ready         (aso_splitter_0_source1_ready),          //               .ready
		.aso_source1_valid         (aso_splitter_0_source1_valid),          //               .valid
		.aso_source1_error         (aso_splitter_0_source1_error),          //               .error
		.aso_source1_startofpacket (aso_splitter_0_source1_startofpacket),  //               .startofpacket
		.aso_source1_endofpacket   (aso_splitter_0_source1_endofpacket),    //               .endofpacket
		.aso_source1_empty         (aso_splitter_0_source1_empty)           //               .empty
	);

	error_adapter2 #(
		.data_width      (32),
		.in_error_width  (6),
		.out_error_width (1),
		.empty_width     (2)
	) error_adapter2_0 (
		.clk                   (clk_clk),                              //       clock_reset.clk
		.reset_n               (~rst_controller_reset_out_reset),      // clock_reset_reset.reset_n
		.asi_in_data           (aso_splitter_0_source0_data),          //                in.data
		.asi_in_ready          (aso_splitter_0_source0_ready),         //                  .ready
		.asi_in_valid          (aso_splitter_0_source0_valid),         //                  .valid
		.asi_in_error          (aso_splitter_0_source0_error),         //                  .error
		.asi_in_startofpacket  (aso_splitter_0_source0_startofpacket), //                  .startofpacket
		.asi_in_endofpacket    (aso_splitter_0_source0_endofpacket),   //                  .endofpacket
		.asi_in_empty          (aso_splitter_0_source0_empty),         //                  .empty
		.aso_out_data          (error_adapter2_0_out_data),            //               out.data
		.aso_out_ready         (error_adapter2_0_out_ready),           //                  .ready
		.aso_out_valid         (error_adapter2_0_out_valid),           //                  .valid
		.aso_out_error         (error_adapter2_0_out_error),           //                  .error
		.aso_out_startofpacket (error_adapter2_0_out_startofpacket),   //                  .startofpacket
		.aso_out_endofpacket   (error_adapter2_0_out_endofpacket),     //                  .endofpacket
		.aso_out_empty         (error_adapter2_0_out_empty)            //                  .empty
	);

	eth_gen #(
		.state_idle       (0),
		.state_dest       (1),
		.state_dest_src   (2),
		.state_src        (3),
		.state_len_seq    (4),
		.state_data       (5),
		.state_transition (6)
	) eth_gen_0 (
		.clk       (clk_clk),                                            //             clock_reset.clk
		.reset     (rst_controller_reset_out_reset),                     //       clock_reset_reset.reset
		.address   (mm_interconnect_0_eth_gen_0_avalon_slave_address),   //            avalon_slave.address
		.write     (mm_interconnect_0_eth_gen_0_avalon_slave_write),     //                        .write
		.read      (mm_interconnect_0_eth_gen_0_avalon_slave_read),      //                        .read
		.writedata (mm_interconnect_0_eth_gen_0_avalon_slave_writedata), //                        .writedata
		.readdata  (mm_interconnect_0_eth_gen_0_avalon_slave_readdata),  //                        .readdata
		.tx_rdy    (eth_gen_0_avalon_streaming_source_ready),            // avalon_streaming_source.ready
		.tx_wren   (eth_gen_0_avalon_streaming_source_valid),            //                        .valid
		.tx_data   (eth_gen_0_avalon_streaming_source_data),             //                        .data
		.tx_sop    (eth_gen_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.tx_eop    (eth_gen_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.tx_mod    (eth_gen_0_avalon_streaming_source_empty),            //                        .empty
		.tx_err    (eth_gen_0_avalon_streaming_source_error)             //                        .error
	);

	eth_mon eth_mon_0 (
		.clk       (clk_clk),                                            //           clock_reset.clk
		.reset     (rst_controller_reset_out_reset),                     //     clock_reset_reset.reset
		.address   (mm_interconnect_0_eth_mon_0_avalon_slave_address),   //          avalon_slave.address
		.write     (mm_interconnect_0_eth_mon_0_avalon_slave_write),     //                      .write
		.read      (mm_interconnect_0_eth_mon_0_avalon_slave_read),      //                      .read
		.writedata (mm_interconnect_0_eth_mon_0_avalon_slave_writedata), //                      .writedata
		.readdata  (mm_interconnect_0_eth_mon_0_avalon_slave_readdata),  //                      .readdata
		.rx_data   (aso_splitter_0_source1_data),                        // avalon_streaming_sink.data
		.rx_dval   (aso_splitter_0_source1_valid),                       //                      .valid
		.rx_sop    (aso_splitter_0_source1_startofpacket),               //                      .startofpacket
		.rx_eop    (aso_splitter_0_source1_endofpacket),                 //                      .endofpacket
		.rx_mod    (aso_splitter_0_source1_empty),                       //                      .empty
		.rx_err    (aso_splitter_0_source1_error),                       //                      .error
		.rx_rdy    (aso_splitter_0_source1_ready)                        //                      .ready
	);

	qsys_top_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	st_mux_2_to_1 st_mux_2_to_1_0 (
		.clk                          (clk_clk),                                                    //       clock_reset.clk
		.reset                        (rst_controller_reset_out_reset),                             // clock_reset_reset.reset
		.avs_control_port_address     (mm_interconnect_0_st_mux_2_to_1_0_control_port_address),     //      control_port.address
		.avs_control_port_read        (mm_interconnect_0_st_mux_2_to_1_0_control_port_read),        //                  .read
		.avs_control_port_readdata    (mm_interconnect_0_st_mux_2_to_1_0_control_port_readdata),    //                  .readdata
		.avs_control_port_write       (mm_interconnect_0_st_mux_2_to_1_0_control_port_write),       //                  .write
		.avs_control_port_writedata   (mm_interconnect_0_st_mux_2_to_1_0_control_port_writedata),   //                  .writedata
		.avs_control_port_waitrequest (mm_interconnect_0_st_mux_2_to_1_0_control_port_waitrequest), //                  .waitrequest
		.asi_sink0_data               (error_adapter2_0_out_data),                                  //             sink0.data
		.asi_sink0_ready              (error_adapter2_0_out_ready),                                 //                  .ready
		.asi_sink0_valid              (error_adapter2_0_out_valid),                                 //                  .valid
		.asi_sink0_error              (error_adapter2_0_out_error),                                 //                  .error
		.asi_sink0_startofpacket      (error_adapter2_0_out_startofpacket),                         //                  .startofpacket
		.asi_sink0_endofpacket        (error_adapter2_0_out_endofpacket),                           //                  .endofpacket
		.asi_sink0_empty              (error_adapter2_0_out_empty),                                 //                  .empty
		.asi_sink1_data               (eth_gen_0_avalon_streaming_source_data),                     //             sink1.data
		.asi_sink1_ready              (eth_gen_0_avalon_streaming_source_ready),                    //                  .ready
		.asi_sink1_valid              (eth_gen_0_avalon_streaming_source_valid),                    //                  .valid
		.asi_sink1_error              (eth_gen_0_avalon_streaming_source_error),                    //                  .error
		.asi_sink1_startofpacket      (eth_gen_0_avalon_streaming_source_startofpacket),            //                  .startofpacket
		.asi_sink1_endofpacket        (eth_gen_0_avalon_streaming_source_endofpacket),              //                  .endofpacket
		.asi_sink1_empty              (eth_gen_0_avalon_streaming_source_empty),                    //                  .empty
		.aso_source_data              (st_mux_2_to_1_0_source_data),                                //            source.data
		.aso_source_ready             (st_mux_2_to_1_0_source_ready),                               //                  .ready
		.aso_source_valid             (st_mux_2_to_1_0_source_valid),                               //                  .valid
		.aso_source_error             (st_mux_2_to_1_0_source_error),                               //                  .error
		.aso_source_startofpacket     (st_mux_2_to_1_0_source_startofpacket),                       //                  .startofpacket
		.aso_source_endofpacket       (st_mux_2_to_1_0_source_endofpacket),                         //                  .endofpacket
		.aso_source_empty             (st_mux_2_to_1_0_source_empty)                                //                  .empty
	);

	qsys_top_triple_speed_ethernet_0 triple_speed_ethernet_0 (
		.clk           (clk_clk),                                                            // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                                     //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_triple_speed_ethernet_0_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_triple_speed_ethernet_0_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_triple_speed_ethernet_0_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_triple_speed_ethernet_0_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_triple_speed_ethernet_0_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_triple_speed_ethernet_0_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (triple_speed_ethernet_0_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (triple_speed_ethernet_0_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (triple_speed_ethernet_0_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (triple_speed_ethernet_0_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (triple_speed_ethernet_0_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (triple_speed_ethernet_0_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (triple_speed_ethernet_0_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (triple_speed_ethernet_0_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (triple_speed_ethernet_0_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (triple_speed_ethernet_0_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                                            //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                                            //     transmit_clock_connection.clk
		.ff_rx_data    (triple_speed_ethernet_0_receive_data),                               //                       receive.data
		.ff_rx_eop     (triple_speed_ethernet_0_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (triple_speed_ethernet_0_receive_error),                              //                              .error
		.ff_rx_mod     (triple_speed_ethernet_0_receive_empty),                              //                              .empty
		.ff_rx_rdy     (triple_speed_ethernet_0_receive_ready),                              //                              .ready
		.ff_rx_sop     (triple_speed_ethernet_0_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (triple_speed_ethernet_0_receive_valid),                              //                              .valid
		.ff_tx_data    (st_mux_2_to_1_0_source_data),                                        //                      transmit.data
		.ff_tx_eop     (st_mux_2_to_1_0_source_endofpacket),                                 //                              .endofpacket
		.ff_tx_err     (st_mux_2_to_1_0_source_error),                                       //                              .error
		.ff_tx_mod     (st_mux_2_to_1_0_source_empty),                                       //                              .empty
		.ff_tx_rdy     (st_mux_2_to_1_0_source_ready),                                       //                              .ready
		.ff_tx_sop     (st_mux_2_to_1_0_source_startofpacket),                               //                              .startofpacket
		.ff_tx_wren    (st_mux_2_to_1_0_source_valid),                                       //                              .valid
		.mdc           (triple_speed_ethernet_0_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (triple_speed_ethernet_0_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (triple_speed_ethernet_0_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (triple_speed_ethernet_0_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.xon_gen       (triple_speed_ethernet_0_mac_misc_connection_xon_gen),                //           mac_misc_connection.xon_gen
		.xoff_gen      (triple_speed_ethernet_0_mac_misc_connection_xoff_gen),               //                              .xoff_gen
		.ff_tx_crc_fwd (triple_speed_ethernet_0_mac_misc_connection_ff_tx_crc_fwd),          //                              .ff_tx_crc_fwd
		.ff_tx_septy   (triple_speed_ethernet_0_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (triple_speed_ethernet_0_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (triple_speed_ethernet_0_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (triple_speed_ethernet_0_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (triple_speed_ethernet_0_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (triple_speed_ethernet_0_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (triple_speed_ethernet_0_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (triple_speed_ethernet_0_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (triple_speed_ethernet_0_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	qsys_top_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                           (clk_clk),                                                            //                                         clk_0_clk.clk
		.eth_mon_0_clock_reset_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // eth_mon_0_clock_reset_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                     //          master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                                 (master_0_master_address),                                            //                                   master_0_master.address
		.master_0_master_waitrequest                             (master_0_master_waitrequest),                                        //                                                  .waitrequest
		.master_0_master_byteenable                              (master_0_master_byteenable),                                         //                                                  .byteenable
		.master_0_master_read                                    (master_0_master_read),                                               //                                                  .read
		.master_0_master_readdata                                (master_0_master_readdata),                                           //                                                  .readdata
		.master_0_master_readdatavalid                           (master_0_master_readdatavalid),                                      //                                                  .readdatavalid
		.master_0_master_write                                   (master_0_master_write),                                              //                                                  .write
		.master_0_master_writedata                               (master_0_master_writedata),                                          //                                                  .writedata
		.eth_gen_0_avalon_slave_address                          (mm_interconnect_0_eth_gen_0_avalon_slave_address),                   //                            eth_gen_0_avalon_slave.address
		.eth_gen_0_avalon_slave_write                            (mm_interconnect_0_eth_gen_0_avalon_slave_write),                     //                                                  .write
		.eth_gen_0_avalon_slave_read                             (mm_interconnect_0_eth_gen_0_avalon_slave_read),                      //                                                  .read
		.eth_gen_0_avalon_slave_readdata                         (mm_interconnect_0_eth_gen_0_avalon_slave_readdata),                  //                                                  .readdata
		.eth_gen_0_avalon_slave_writedata                        (mm_interconnect_0_eth_gen_0_avalon_slave_writedata),                 //                                                  .writedata
		.eth_mon_0_avalon_slave_address                          (mm_interconnect_0_eth_mon_0_avalon_slave_address),                   //                            eth_mon_0_avalon_slave.address
		.eth_mon_0_avalon_slave_write                            (mm_interconnect_0_eth_mon_0_avalon_slave_write),                     //                                                  .write
		.eth_mon_0_avalon_slave_read                             (mm_interconnect_0_eth_mon_0_avalon_slave_read),                      //                                                  .read
		.eth_mon_0_avalon_slave_readdata                         (mm_interconnect_0_eth_mon_0_avalon_slave_readdata),                  //                                                  .readdata
		.eth_mon_0_avalon_slave_writedata                        (mm_interconnect_0_eth_mon_0_avalon_slave_writedata),                 //                                                  .writedata
		.st_mux_2_to_1_0_control_port_address                    (mm_interconnect_0_st_mux_2_to_1_0_control_port_address),             //                      st_mux_2_to_1_0_control_port.address
		.st_mux_2_to_1_0_control_port_write                      (mm_interconnect_0_st_mux_2_to_1_0_control_port_write),               //                                                  .write
		.st_mux_2_to_1_0_control_port_read                       (mm_interconnect_0_st_mux_2_to_1_0_control_port_read),                //                                                  .read
		.st_mux_2_to_1_0_control_port_readdata                   (mm_interconnect_0_st_mux_2_to_1_0_control_port_readdata),            //                                                  .readdata
		.st_mux_2_to_1_0_control_port_writedata                  (mm_interconnect_0_st_mux_2_to_1_0_control_port_writedata),           //                                                  .writedata
		.st_mux_2_to_1_0_control_port_waitrequest                (mm_interconnect_0_st_mux_2_to_1_0_control_port_waitrequest),         //                                                  .waitrequest
		.triple_speed_ethernet_0_control_port_address            (mm_interconnect_0_triple_speed_ethernet_0_control_port_address),     //              triple_speed_ethernet_0_control_port.address
		.triple_speed_ethernet_0_control_port_write              (mm_interconnect_0_triple_speed_ethernet_0_control_port_write),       //                                                  .write
		.triple_speed_ethernet_0_control_port_read               (mm_interconnect_0_triple_speed_ethernet_0_control_port_read),        //                                                  .read
		.triple_speed_ethernet_0_control_port_readdata           (mm_interconnect_0_triple_speed_ethernet_0_control_port_readdata),    //                                                  .readdata
		.triple_speed_ethernet_0_control_port_writedata          (mm_interconnect_0_triple_speed_ethernet_0_control_port_writedata),   //                                                  .writedata
		.triple_speed_ethernet_0_control_port_waitrequest        (mm_interconnect_0_triple_speed_ethernet_0_control_port_waitrequest)  //                                                  .waitrequest
	);

	qsys_top_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                // in_rst_0.reset
		.in_0_data           (triple_speed_ethernet_0_receive_data),          //     in_0.data
		.in_0_valid          (triple_speed_ethernet_0_receive_valid),         //         .valid
		.in_0_ready          (triple_speed_ethernet_0_receive_ready),         //         .ready
		.in_0_startofpacket  (triple_speed_ethernet_0_receive_startofpacket), //         .startofpacket
		.in_0_endofpacket    (triple_speed_ethernet_0_receive_endofpacket),   //         .endofpacket
		.in_0_empty          (triple_speed_ethernet_0_receive_empty),         //         .empty
		.in_0_error          (triple_speed_ethernet_0_receive_error),         //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),                  //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                 //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                 //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),         //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),           //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),                 //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)                  //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule

// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H:4]0UL+G%6A.UKC@4I^X+DL9N5V=5BUBR>/G4/.K-'4#*&QD9I :1   
HG:_ZP7V/7;V%O6 L)&8U@.1=T*(A%4U#9>MJ<N? G_]Z-!!8P8O.B   
H(0,BGM7?[Y5.IPDEB&SN9%W(#PJ3TE0W_:_<1?WTJRQ^IJ4*^:K?2   
H\1O$&*41N/ +ON"=L>)ITZA-.E<A+"K8OBI(O9-[A8X<LIN63O#2]P  
HWT%2*!B/6MRI;59;C,7=DB"XZE30<JHT,[2S?JG+!6-#0EC!9(1OC   
`pragma protect encoding=(enctype="uuencode",bytes=4896        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@D:"TD.&1(I"Y)"@[P\$4%J&[:!6%2NG8D)*?%)]%IZ8 
@N&X0),KQ_A<"Z^F[,\/S=C8WV_2A V88TB%IUW8G54  
@<B4E!<Z$POK2T8D-Y4PES'N_>!PEK$;? U\Q>H:X=A  
@!N9'(+OB6KYXX99?>1DB%.Z;U_&3MKQ!C]G2"5I'(DT 
@&5]:)*A(SNGNPO1C9E@]5EI)3CN>NG0@CY50=YST6M  
@$W':J 4QR8M-UD$M(HB,8R$4!:N&E5C&)>D A#,A=;X 
@B7ZVRCW:9X^6D;!,8JX L!R>IG%51[B1\9 +,&T'A7@ 
@Y>IWLMQF-CPNQ4D1A5B5 PNV:)U$I)M2ITHQ NE_T>\ 
@%N1@(1HJ]$##K-1H/AF>'CC:L<C](\J-$0.KQLZ<J&P 
@-?E-U@N!4^%C,:?'8<S7H#$\ '<Q]"@F[J33,JZ[Y<( 
@$F:3ZQ;J3_?WG<:2RXI:'>A=C9:>)-DXA](O)5$$340 
@Z\_@5V,UITM607O$B'H;#+$26+FM6V)]M["+@Y1=, \ 
@0%ZXV'@C]G!N]>\YV'R[%"7[(!WOKHIZ@ E$4.;#+90 
@I2"/G)B6T@3 T>LG"01;.6?1V'Q@F:,U+OU@*)OOD^P 
@RD*/K\3Y11F1F]<Q:[8XL,!>![-DE_BGVS,,]()'Z)8 
@J@0%&F]G*#H+YKP@;I;G6\6:FA!X<\%0'\Y+U19,,4\ 
@>[!$3A$-NRP#/F]#O0T]PM]FPU8#/;Y5JE42$HP(RQ\ 
@H:H[]<OF\TU("ANJKF:1ZD(4X;<#*1Y1JWN()2I'?YD 
@D,\7[ ?JV=<!O)L\V(1R_(U>(UTDCXIBE$.WN'4 :?D 
@H1A#H-T0S/9K%XFO31/"TAG&,Y)_:/?M=& 6J-NA,U, 
@1#"[MKG+JGD*%5XY>TXW$I!;_UKOS^"PEB^G5,-!5FT 
@O_OZ(<91P2.]#+D^)3&*W/)NE00B<86-"[P"F9F<@Q< 
@>G1!@=(NN9T6G!ZI;N%Q?93MP6OJ5?0N(?8G-0*B-YP 
@]P:XOI0J^>PQV?$-.9%V5Q!MY=R!"NQVQE*/PO81UI@ 
@^? ^O\L?6V2RB?VA^"RW62,B8 %^4K*=-M8)@EQ"%H\ 
@:%'[K<,2.3L0 CQ^3='M5C!>>F477=QXUTZ$6+'EEM( 
@&TGS4!ZA&I,EW#77T>#H^W 84+<MQP>B@-)9,[?3XWP 
@WV'+\\"JKMJ=9(6AW!C+KAZ&U^<6+*M_@NN\2^0H)>4 
@OK%4$:OB<0L:YA>M454A&VJR?L)Z5U8K/(8,9(Q8=60 
@EZ$]#YS$JJ5 72</W=])8W,F9QA%S[$N:>*3VX4\#F8 
@\Z1TFQ!!YY!X*#2+ ^@\0T$;ZS%_"\ 3A7$$0-P!'/P 
@/^ 4<P=.^31J,,0YM]ZG3JK2(72'C!>/K!Z_'+_[9<8 
@#2=I1T9.+)5"CBAD;1,19,_+Q';"\JD*-J-37P_YND0 
@55QPK,&I=@12FV4P_NBG94"VU/YP&1TE25U0F4RI[A( 
@7DH>E@'VX)#N+1)6T&/<V?\LDR ]*+,;*QQ#YE<CKN( 
@@5F?L@6< "@7"6%-=0P:FA%)-@ (47]S[\0W-@+H8IT 
@]B=$_]N&7W6ARV(&9,Q_W:)K(FA:><RD2Y![K?+CH;0 
@!BGV"C,=O/GVR7A:&T\RS-*+0""#D^.ZT?];.95L@($ 
@N;N *6L<1(S^RZB&Z "*+-,F7>0158H9DZ)^$6L=>H  
@N'A0S'O5^ZP'UW0O=/'B-AH;N&BM-DY$X7HL6 L>=4P 
@K::M>4T6DY(S: Z[UPMEXB16>3;6R<0MO0]TL.%_5^  
@X6OQ<WIS<)VB)>V<=F"U]L(0B.:7S(!53PH#>6/PCV@ 
@"EY%;=-QZEN*9?H-KZ$[JHKR\\7U"PO1M.C%F8B:M,X 
@D?L)*$-NG)PUE;IZF9@+NHH"(;/[\2'?X</^!IB.+FP 
@2DQO_W /?19)AP^=_S<O(&U\[%G)"/0,X>C6*HG?<S, 
@[9Y=RYID)>.ZU:[3A"W6Q$V(<Z/T*LD3,6[Y"1P_XRD 
@5@9?1R]5L,#H,(L*@B0<Q4@%1OD/_B^^2!UX,;7KOGH 
@+&M=<U(&51?M]%^V3J@LD8UI_'XIB$VQ[<EB,:SC 4( 
@@ZB$G9@(&#[@XY>YD-TF?)5WP>F$W$BVLLLL/8=>B6, 
@EXX/@SJR5JKLEX[5L:SI!P1?&39/L*S9]7#17;PO228 
@EA!!(<GB<5-<Q"HS/_ 6)@!$U:PG(O73ZD5!$1R"UNP 
@DZWD'Q'LV\YBB"I*&>Q91"C(?NOWS205:ZG7:GIGJ[( 
@:&KU*X&>!S<-.T>Q=/9Q?HN>Y'I4Q?T7Q0[^_F>^BLT 
@_5?T4?7=V=4'>FER[=.!FO<GR2+IL5@#JJ1&JUL*,1$ 
@E#4FX@/2R6@H5G85_LH$S#QX+'IG$Y+C\B6F_U$<)44 
@_K/Q^D<)BN5:[V075J\_#7S"52;7_Q4U/?[EN!>=60@ 
@KC+3@=XATH8ZM->45ZU4"X7PW-'?B9">N:,)U%GA6JL 
@_W'66Z+/2F\>:64"P!#1:7OU G(F"2XU(.:3O6']@PL 
@77SWGL-TP\'='5.Z'HE=91Q(>38LTC?W+?#';+S;SW( 
@LWX_-^/*)).Q=*=F+NX1R[G,+W6QV<,%UZS7-\@J4\P 
@=.&CH_QI@B$H3E]6R'1;U8CD68_ X8H?V(MHEJ0;2K4 
@"?,S\Q(/*Y2_GSR"/G82[&]/*2>-V9.]/=5?QQ(_GF4 
@W<E[H0ZN>W6<YF;F5Q!0E,^4!]QI/P(^9_5=9/C__-4 
@+LQC/2T( ICZ9 0_7:0'E!1Y4IE*3M!C1<DY'P=T+XX 
@P75U.#^LV34+(R@2%,8/[H;!:>N+.0K*3T0A!H8[>&P 
@:Q-ZMU=,!NF\GB,-QTA_1B9ZT34ZD8D^#PB3<^&((70 
@/U":D<7E14#B@"3D!+J3\A-V'';$XN/B3-[B$ !(%<< 
@*>4@([LM Z!N0F//[F84X;ZPX(!%BS]L?@X;J6[4.58 
@Z[9@W-,Q;J&6%38E1J-RY'^<$434Y2#>=6OF5[7Z)W< 
@&5!@5LJBGZ+ !FSHBR<"/;V$M\A]"S+T:?.,O1^$\T, 
@-71;^H*"DX<V?GAESR@@:$Z(LX";1D'U7ME])=I5F<X 
@ U,.$V>/NTO$&%),#353]RJ!-XGA5L9Z0N9J0BC"$^D 
@>_@EV7=QCY.PE,'?G%0J'1T<5>7\(D\+(\LE GCI!ZH 
@V"YYZD[?ZE8!_'-[%'\".4'@Z1Y7N<6\;ABFR@"/5$H 
@I$N_5B1/Z@ W/46J+EKHLX3\:'",S$KK&!$D,V+1YI( 
@%75<*])P4;&;2G:#@LQQ.F-AR;;J(.IW\$[TVGK/UO0 
@FV@<'_KO\+M&.2!W1$]0-U6RWRS>KFH F4#EUJYC6M8 
@X7Y(('@DK5$UDJ]/)D5Q6$9QZJ:XPT2JK/.7S&L>O]0 
@$>>/])M5%S91L-Z;^)P:471&$*E^'A<89>>=&-M*:O0 
@Q>B P&,7) $^D,5A004/=1[I0$F?D%HO@; %!>F.(U@ 
@W&XG!'?2(M]-_7Q0WNFG&OG^(+*PVKWEG"&17!NA+K( 
@HX"G F,Z?87%O$--#3>G/]>^DLQVCRC6P9S77;3+L7$ 
@KJ/QWXI.9O.I7J$G@T$ U*DJU6Q6,J:QY.^2O]EC'*8 
@#\&9K-TNF+63O*X495N2_81+*F>!LPG*DU6KISF3S,8 
@J!]1D&2;*Q?'1+ 0\$^>!.K P$.JJ2B8(Z@&WK]*U-X 
@PKFEUMJ5_.[@% ),$Y%X4:,*+%Z_'=[KE(L>&IW !TH 
@\4P9QI1$"CTS?_NF65:Q!J4O7@E^Q<TAVW@S2;=67;@ 
@T2%CZ"X^5S&(XH=L[_,*.4&O#A)8)"\,X:EJL_CZVY$ 
@IZ(_A63,_(5F$4 ):W>3?T@,D\NX;;X[[J$&&1J945, 
@I\'HD7E^E!F8P4C(PB&N2-P!$C!_JR><NX-ZV^T;P!( 
@<Y%EY^\C')H"[0TG)UEX^OZ]T[I3E#FV7YV)YUOQ0NT 
@R67G)GFG<K:M:NT<I(/Z*W2L6#YG"7,!IBK:EZ1K2HT 
@3^S*#TB7I]*QKY*2(6N0(B!QQ5N^*.E6]9L6_11"8]P 
@DN"KX;]744@7)8($'O\KXARI:!/.L5S<.D_LSSQ,Z'P 
@UQ7"YZ#B""2; %?Y2E W/^'3.HN@YD"(4I+)J,A(\2  
@[+UHJH64^V,J+(-H08F]NZ'8L1,%10Y0?5/ +^@O<$L 
@$\)Q?VKU>AP.&%YS-\@<?]D'1MR[,N5@#'#JEFT!JH4 
@EO.6> .<(8(_9TB4:6$ 7/]&4>6V^<J^QT%+T7^V\1@ 
@+1]'H*1120D@Q^ARI?L*EW^V%"C30'Y:G(C@ OR#_+$ 
@?T.Z3:FZ2]^?>QDEI(YTD+:(<S2SKI?J*I>[QHT3;J@ 
@&MSIVQ C9<[[?<HVA6N C*,I:E$.!E720\CEQ !?%M< 
@43YMG,?GAGS9$T4_Z:M&AN")R3,&5@;W^4E,9+0B!KX 
@6U"QUXHSZ!".5R1DD:$J]A _;_,Y!^V2HENEM?I<<4< 
@IRENTX3>E4-=P[_![?I%J>7'(J2P@Q4T8?+NKNKVTV8 
@.0VZ02:!JZQDRX'NB?<: ,[< W)F-EPBQGL%C[0:R(L 
@]G0"2!JUZ]+8]T_&#W.P?XBV>&06>,718E)CN3)\ TP 
@5V^H]R* S&/WQ,@8H)J5'.&829HI63@3-#BC;X2QN70 
@B3E.S4'P*G@U3<W%2^]5>Y]5U1>/[I6&0*^X<G*W35, 
@CF%X4*\X'S=6\41G;;;=X2\^QR==,K@>"W)YX]]*G,, 
@/@[2L55#C&MU?>]LB6VE%A/;@I"J?GUD5LCT55DYPE4 
@^XCIY_WZ0"AO(=>U>F#KYCW9;2EX1)D=:I-22,UZ *8 
@3X)7YG&3,*S? 18</<XBFB)@1:]_(0PB7YB*F]8%X*( 
@9F 4\6/V*XP9/\D:MG;SV.5ACW"[+74.[IE%/H%1XN8 
@M894!.-A]N""):@"U:2I'-$6\T-#N;F/I ;*(!U@\8( 
@JSR(K3-[1.P7<)FW\*![$4]LW-6>DTC=G0=^YN:@@"X 
@9;B5C157:8M>\6H$I/W'>W9D=A7A5G:',;RG,#G<Z?\ 
@]D(?!Y]CJ)#G](OKVM, \&%%+:TQEOP/!E/S!F^U4QH 
@SYXBL!HJ8OZK#1B-78&'T,BY5.N&<#]$%Y1+*R,=?8T 
@@_UU'"9O03A%GF\TIV=\QDR3 8"+9,+C<TU90O(G"^X 
@G565PLDFNQF"!@)M*KDKJ=E;IVBSHBOK938W'%H%R%  
@#T!7P8PW7_JL))D-N09>1<H"_"XJ&>K@]7_8+>)S_>$ 
@M\9[RG/_=65T,4'G!!(%.2^Z>>K!LQYQ^B$<0$!XM^$ 
@Y!.,+8)\BWVY3J#9";\F10T-D_-\\PI[&%!U*AEIUO@ 
@E0^76;_Z,TUAC0I,+X$2#@6'4[:='Q<8Y+N^^[S(T)\ 
@2PHB]@=GU] U;OG"):(%8K])&VD[@%V+SK(Y5:M^&.H 
@;C&M(IHU#X[5%V,>]31.<27^E4<[)>O@'WQG9<H<!+@ 
@W5PX@25&Q4^M:Y?R&9V%GXPYBD"*A1TJ%G?E=MR*>^  
@9V@50^_"6Y'9M,38H98J(:8Y*[&Y;]>2^UU9$%F%'DD 
@:X#?6&ZIR_BY3B"N2D774%6?F<%LK><'-Y$>Z(; %=T 
@N Y?S-5+[2 ?9BZBRA!Z8/,3ZXM5I8.L6ANZH.0+&_, 
@%D#D]BS!+!^P9JD_K)><O6?UA.JYD<<LN[4BXS?XQ.0 
@:?C=UMLH'#3=2(9#.*BIE_TQJXMC!XW[&BZJ:AXU#S< 
@.K@H;O!-X;-P7">41[X X-P"7U]:H)A$NZ<Y/O%>%_D 
@])B=FG&E'X6=(:PXQJW39ZS+F_R=*ZWH$>S5HS-YR?\ 
@[G!_&_=.DAI//(_[87-4C:8;9+6-0$'-;*(?G)0SL28 
@E8'SD>K_Z-N-5<!!S'-'ZOEZE]AR5HR L(Q>N_)UGG$ 
@9"F:D05J#@S^ZW##?U1 =)E?0]/+GI'"<+E!IWS:)74 
@=5+92C,N24W4G(8,7/;=OJK(_Z4%SA6>N?)J]_C$N)P 
@T$M;KX MEA  ##E+@$>&D/%_#XDQB?)5 6^@QW.B2O@ 
@Y;!_?2]BZ-*A<AQ^FJ]Z#WYANK'N9:A:96'O+56I218 
@3LV$1ELW504W;RO"!+WK&!![2WF0;<ISO62<KC\2W\@ 
@K0FZ=:Q9%X@53LRZ3[Q?A_I45J0853^CA(B(R?Y[N4< 
@4*.SPV&]WFH^[H'0B GY;A_70HSHCM47AB8+'680UU( 
@UTYH>,97(L]Y;50&$CARC4G K%7, PM1&B3^;QR5DK$ 
@9K5Z*]H@0X]&$)!"8!K6J+^A50Y>VW0(&< _Q4P\9P8 
@MELL6Z4F*4(*,27%8);"E.VL,[S6KUZ)@;=L.JU% 3L 
@MM]'E,3$'*RN>3N%<*M>THH83#@A4HEQ<[SBJYO$YE< 
@$WQ*K&RF]G]+ :3G;I1L,,&6"8A9TRIP!AL@U?N8=AD 
@L-YEFUUFM)D-;"'LKJ5(]8($)QJ<-^7>/Y>3/1,A-,D 
@?$^) ^\,KN;_#J09BC]_5V)+C>NBZ@%1']S?E(^,?]T 
@_$Y8^#B*FN0V.P:&4U$&G*%6 _O05PBO6,%^:!-/18@ 
@9YF&WWL3S\IOZ!Z\5+WTUHV9UJV:U<;YH%,;#+:GVE( 
0,=EY:!B89G?\/=?<&#0-2   
0L;6\@+?JB_U& HA>]>!*L0  
`pragma protect end_protected

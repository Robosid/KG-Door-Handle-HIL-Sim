// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
h/6U6t+EQm0xfIeySrz3PAzWG60rvT+ADrdgZ3/rLBfNYCHW9ByeeWYemFidCbNt+OM/p3i8f5ky
rOZeUE9Pd2yRtk+DCOjkFuBB5HhkcaebU6C+9dN6SrK3my4SoUSMGLLaKbzm4Z2Ww0ygIaCAgvJg
8fdYsbSaZ1l90gJSaBafr+XNbUgrPKinT57/jS2/nUjQqjFCzJx00P2+k5vCBJlGatJe+bH4TBUo
Zo7yyPcJiHoL1/aEGqmA/DFQp7ObDGqhW9/uVAk9D8kYzQt6hnr2d74lvCoNR65R2de05obvzgEm
mowkRCNt/sL2gO6DSTAyNZ9cmY1wgqXUNoHyLw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5104)
brwr70J+zo102ya0E8QIPXjFIBHySwBuQ/yEXM7gp5kC7s7PF333kyMlnX3B8fcGieyDp/+n4aSn
PbI4SZo2evfnBH2ONP2vRAvwcHQmWbGSlVaVAkCZs/1W1/7oC0oLegNn+HoCu6kHbYyi9USkA2oh
QLBA+CJbg9j6tkMvTQdgKLkjyrZMoWN9J6J0ft7PBwQKIm7RqdCJUkZyLZf26rJG29MLGW1pDH/e
W0xoyRZdtPjk3tS4ZgK9FtgM1zgE0xCfuk5XSuZ+Kc+IQ561uhnnVm8Gi6DnAxN4Cn/DWy2jRy2k
gIy3nHMmrwCBH5uj1H0yBo5xnHak5vobiS4vWKjHOQpL0oGmHfSb0dWQstapRp2eT9XaDSW4bSh7
BkXSMqO42bUV9pxyLsX8NYCNUnCY1qOY4sbRDkMR8kfT7jbs4w38Os3R+1wmHQ0E9eupuC0bW6/2
jgXrWQ6a+7k5xZz9EVTC1u/HdXsyuEwDoByo/yi21x5dyS0BVstsACjCykzYV6k2WRAal6hH9EI/
pNI5QyC84fi4O5Z7GM4S8PnkrHZ/sCLz36RWOYLqQROPMFQIBrx+0u8AMATJzxKSUzPMGi4taXhC
32vTGzoIUMa5L96OeRTv6MP+vOuom0dULX9hA31XkQFYmdoFQhicfGDANEuPg72GB8bRchu+LovX
PqjJM0r0gtbdEqnAxDANn9d9dEfOdvqqM2NUqTP8DH6+gTiB0GRplZeaWrJJI4VNCo6v3CIOx4K7
AHDdOeh9SeE58WnMg6vYc5vch0mcA8/Qeu5ve57E3lUeyjgO19EITCP6Tbm9bWgjSfSInwGFR1XJ
bGNo1GFXmLXw/PfYcHxIYEqcuwSzcs2KP/1L1u/JbrsyqsuMTHa0b071fc8YC29XfHgcYUHSuPmq
ow/FJvK+Q0tIo/BpTR4AHVmIqxuaXuUOsEEHrqkT0J1RB6s8AAmRoJfONCeQp5RSCkLHOt/BlVJu
A04baX+U4d3UpamCtbutE58dO15eNqjFOHk5JvLPMF1P85lRgXJVySHckzqs5VnuM70bZm2dqeaN
U+1uX4/QYz01M0YO8ip0eE73Fu2NOGe5bp33ayCI0KyETR5NfvLgznrWDVfsWChUrQ/nEGBiTZ9P
zecTJmo0X4pL+Ihblpvu0Nsqrh52hbEAtUsZyIiqIY0pi2OjjZ48pIKoXAWKgQp6OuFAlmNU0vvE
lL3ixx7YPgyI8WxBZaz/fsnQtBtnEBhXED7QrK+FXw0BSAYrCMi97MIH+QRMXiWeh9VQhVT2rK0u
vxad/JxRUZKrgQANPnHOaYVLRK8s9jyriFg8LQbducMoo9IKbZXUt3NkJndZ0AF+U/acIjAfgHNw
Pl2fy4KysDLDgv6M65U08FsUs74VhR/QZFLqB1Ef6rhwkd78DJ90IPIYmlTdZ1GrZsb5QdbQepGi
b6GU2CNSbXtBKw6DOPHAngtNND+xHZqGtmxsIo54HzTEPwOBmYh+8vu+OcbvT0xp8npz1l20+maE
YgS9T/Keepf362ElnIfM4vo3I2FcXVG+IFXmnH9vVXx3BlvhzPRdjJellpikiDHN4UFubVJGPvTV
M0FG5ZNnsQMBNvnS69L6dMDL8oOcHHt4BtnRc6wzv/GJKI64aI7ivwIc+uzrnFI4D3rxTSoHGmzF
d/HuGpoMPtnmrJimbnMmZKZ09l6nnn0jMOlaQ/QT4Im3z6ors6z5choyAMI5NBiPZuvDDmaTLO1n
7gNhwpNzy+WoAR98cvkLU7piA0DbLFYlSGDtYvBlkyniN09Kpow4YEJJylrGX3L3OmkF/izJJzAp
fNhjxThKUGqP974qZc4SkC1DqKX7u+zvD5ZlbFJrWjqNBYGvRD7+V5pRtx8yYLbkAlGNm0uN6LBH
jrhU3EQZej3Ik84KgEp2R9bYgC7mt/fNF6bbriZsDn96unb4H1zuecfnpH5jR6z9PGhB2JFbsrJW
6BrvuuznypE9UtQXLD6nGAdTicCyXDeSFv+I5da5PMQ8p6HmWH8nPJ7XAIIqRzsb4AxiRMWdyr3P
TMmvjT55mqYiNbjnO8J58GUV4lAju/q80rRiXMgYOmjgD95jgKMYAn4jVZ+/F0GbUxsMqWWieC77
vouCazyXOx44ZoBBOZWyIeWsgnD8aEvBrs2hoKEuehFkK8t11pCywn+E+6rAAl8SLaCNVrkzoCJj
x73wqMZSU8oG5wJj9tZqciFdQNTqkUreUE8VMbiluOAGjts5T0yiKjzQSC5BwMCG1PISrkWUFKca
aBjUNwW6JqwuySlxCHr3mvMUALL4jNW0ZHq5QJg1KaBijl+7M/vsBa7cG2dBS6wf7cOL2aS5TJCE
599CvyDlGuybDyzFzkV3UhrplQgIQ2s6jYyXVMbjII+2DZQPUr0pOBjT/5Pwqwvoxx1w/l975HNB
gxL5XYLN9JvaCv+tzaePi79xYF1/2qB6taxKYpyhGEkm0GBFVL1s+fVhpgGCBzfDdLPU6Iqqtu0M
32mRaqkHD4SBbGVl7W3L35CcR/lzlQCF+cWs82wMZiOHrsk+qYOqBGJJgmP7Xqcsxbpdhg3OjhWB
ObXTjXB8WnR5sT4zuyljjyNAS6TNqrZGie597FX9Ixe4dCrZNg7qbvb3ZwXcrMxggp8fOEsq4o6b
RMwSabXMrGE5qIgjIFOxNOtX1GXRuRo249XgXAhPK1jHKnY7rntpHQi8zJkIqr+AsqnXGEI/XX4z
grSkcLAzQ6nejIWwo0Rt9E49nvZcncBVPlEHXyn/k6ijrvoyuJoZyxOsHMqH5AO0Io4sz2Vy5NeF
1UwM62yTzOwngUyYdKut8BnwZEfa1YBeud57DuqGAzTlM2NrCYH7ghNfGv+ZkICc2D/P4y7jpcI0
tQZeiGZCwJovYTmBskFES7H36tEcpDsUpC8uNzbJZdSAgSeNZI1pMJTSBcsfozycX2KF+kK8afE8
coIOhHeFoeAxRUDSWQ1ljnaVlBFnduGNfgjyPMR1rAw4xku9zAKrFutcwSwfynF45ycvAzAgw/rv
V1226JZdKgfDzl7ig7N+ZOwCIM+jV4SANYRR25FfOHpsh/BRvXsNwEBMwogvy3A5perK2dHx7sFj
gog6UhV5SRO5WipqVKIbZl8Sw8s9ymewEWdFfiHQMqv2X/rqt30CaI2uiqCiG3spCe5Xjk4EjShc
3ggses21t0EKzs0f8TcRUQMnN7TLO1LdPKtp1ottd1+Js0Q60nxlUzNabfOeu1EW0hGiYMiHtpef
dmUq7FjTjUswLS4Cj0njgm/G4JbEkkWGWlLIwnXSV4Nx2uNvwa/F0A17acHYthnQjnn5PfyRbYf8
KKAmPV1NqCurS+dAWqYGkV5yUHVLjRTVY3KpHkQA2ZYIeejnSdLDqPe/XUxLnApoMcuMAyV7PsSO
FxQTum7EkjWSA7PSUSDqOxyC1MCnJdWu8p/bSPsH68U3rb1eOdHD6WQVT/EQQdhrbiqvUQI+wK60
+Wx2fxx9uI6JCNlFWVpbKT11UfyOTSOcrYR4QyvmsrTInYqvcPaKixOBK13tAg8RrF1uwGHY03ih
EqJLx1VlliwbvZpa8j6lX9NRqeLkXo/re4ptwsV5hCr1uEsmkKIN7O542bLXM2OITMNulwJXKwd3
wgZ0hCpecziFNeTb3y536BQpkzfli7GatLROZ7pboyBl/+FcQqF2z8utKI9M+G0HkavPO9Zg1Xxv
022MXlgLpcg34udAUBiTfOdSKJ81JN5PU75bKTXqzIwZikMbOy1/KNUfysRObyyu7WkDo58nu6ub
JcMJl3wmWhSrtOVFNkAlPtIpay+0RAEfnBc7K4ZVWGAwOjp+HmfwSiUXlx0FdqADzdfMTa+bh9mF
dVszqM6W+3FJVPC2DDs8LPHnbAUrKv3E0TabvpEYMeVZ1MaUsJcQK8ISNKojOS/VIzxKW8Ay9iXz
Edzd/Vt26UapqYdXRJvBjPO0R7ROXIr47LsFMlqhrdXz+r/3O6KrcGTye1hLpkuIAyvzMWDUDg8w
Q1VpDdGhWlodnkNEa/dP9Obq1uuTih+SNMEy3B8CskBqFzSplsWAILI0u+f24y4FM8GXDESn0QZT
LUxQGNSxV0vG7Rf7pmGGoksI3B06eQ/cEaZVYRHf5CHbYMzNL4XqmQxexFt0L+gFEOQlymOfDBfZ
pmd+NVW6MsPugQyFq2J3nT7/aVc8LJTqgS/kANlpyD3VTKmNo10hyBKhSJMIu7/CRVVtq1kSrcTj
vHlIfLA/cGrfBu7/cSwqWY/I5jlCKE/DMCqyvKUn26+BG4H449XtJ3FHmFTdgJVOZpuvvmIrbpPr
eoFuKo6o7IfTiE3wTb8oHcNKsHoCivxbgjq6nSMrj3Xe1YuVVfZ97ds8gJQKyRCc32dDpX8olp0G
HoNiM6ZEvY71cuVXNDCEAD1XH7Xs7saq4XbsI6C5wXXPb8qfw8JsWYZcMuavPvVLDqozpNHp90/4
2mQpuyi3nQWJsg5KoVlbiffemgI/tRrfgsFrd3KBM2ogS5VUMiDDOD0pMZoo/vUGxoACQupZw0EG
pBKvmOOqwlLiw15l/j3DvhyxjNm+RqqpW7tdVQMBHkn93H4oyOe/xTDoqnBug4h00XMoLNXu08W7
Dqs8ccLJ6rMQP3/ZGbqw5DKPDkQ+TdAcqGQ9Tmrl+AOeFk9BhC9jWbIJcFfdGpy27lKBhP9LLHOo
15Mzf2hGwrg1ma9l8682MMF+rLt/wG3/dM28HSRDdFoCg+JiE3s5ll3mgTphLk2UNImgT/Zh1zKn
+pc3mi2SxJ4/SzchNHcSaEZsS33ZAeKlA4qhW30EcBOFsi5XVJABvikgj5Z3IxCF3YrUDjlf5Trv
w7MHAEN4V57fpzvvdoRsSyLIHbwQGUeLx+rvzM1B2+BGRc8ZIKxtULNjeE/NG+D+B/369Pnr6Mxo
oXGW5jTgt2k7tbe1mXsI7+UHVr/kkcMW/GnsImzxxuS+A1JmeQlu1csWzsU7K/vBtNu9lQ92TKuT
z/dwybWaSJ7uXTuEUSDKQwC4mwbsOvyGr9K3pijY70RUgdx1DWPKwq5NO0PBfZ1cW1R5v+mqVnvE
DjetmuRFB4cijC+WH8zW4Ci9u/UZ6vHA2KeJ1YJOC4fLk18qvI8ZRK5gNZXpFnH43CmEDhj+7SML
KQcnUdFBQGkAsZOUjI9llj3y9u0Dh2BvWoEctHe+Z+0pWT1AbscBgu4NLFaP0TmPCQL0u/3rUvwO
NXpwHze/SXD++PZ8aTA+076HGqT1W6H4SHdPDnXqKD+GWMqRiQmkUi2TTNqhrdbJ5ulP/XyK1yvv
gN7NId/48iaWSy86zKiWyVZQXW4tecstsbUHfCrzlsoKCvVP+zjJWUkQPdg4OHvyi68fZ7lLqytV
q+o81opKU8qX/re5sCR6kZ1rW+X6qBSimWH5seCY1Dw/Zim5jxlt34G00MFbt7p8/UC0P675NgEn
JyBWDaKI6M+KW/fIMi/1XSOfN016cecfLFhFuag09jIQYdijgKb4653T82cE/GiMGlgiYAaF+3by
PZW+91MdmJAygjspIIpkCqyUuze+Obnyl3ULnzSzYeR92QbJsGFjihtJOEecHID6CF1FJ3mVk8V5
p9v2nqwra3Y2MNgt1XFjtdR+jIxNfl329b2HgbzMDiSu/rDNgwp+Y7vPM4L6fsKjkOSqeQHRX76b
b19wNgRxXv3uMv44gcwNCXbYmGrYtkydmrPJ4he1HN2BUxucPrH2mT3STVs+FpNLeEyT3cvG5eQ/
iEHAXbbWNU2bcRGOsVS7dyk7uIyv4GSE78QmP1UfzE1LMVUAD8qRnFyaI9pTgCaMOGmfL4hf9Z/k
iI9GB571CuzT32GCnORnGbL/hkwRu5xQEJhygewCkRqpgaEGgMOnDZHVGyBVERIMn5lGxTHttYZk
bjVE5A17keDqzweSrQsyjLK+J7osFqDsshCckULB7eGiukGi1Ml0S6PIhHn8zYTI1WdmZkR8/tSO
QPAIPtex2C7x6uZY418KUs0pdODpDqPAEgzr/nzhWSwa477/ZFWxMuIAUHP5uKebtWYZywLMOuaR
Tn6+02Ell/MWa0GMXF99tVVg2riMdRlzYvGIr6Ol/hhdu9oFvZFpdETdS7FN1NxNkOUsJAZ5Y1qG
pbekyow7oskcY1/Q/++zReeaDqnR1YD+ii+VVeojwwYj/cACaDUgqroJngNW+uHohaB2jNY8RbWa
zrrb+uFmWyAO3mYlElUF9g0mBq3Qjf0dJIFV7V8RtYwCVRt3hSP086zA5hAWg4wywLoWCsbK4JnH
SnYLpulDV6VAlLnOxutbJMzLHry6gMy3HSZROX67c9AyngQIgijeAIcqQXaVOhqhmKCCX7d/s+Qm
NMdMD4CRtYTNPLjyFFz4KUcGka7BoAzYxBL1/2ehjE+j4VtQDr9D20R7Zx2ewZOlvhP9efEPgpgI
1dUg1W970gVHxso+kIBHAVxuwyRe+lmEBBXdk6O4kCi0+mvAhp5XpH2niYxXS8Ifk38jaKhBFTz3
8fYk4byvrxfQgNXm3iPQ20OU5q3Zqprl+zErkakO7YkhgGdLYd/oNN9qJ2ySHj37TrQLMa5XNtE1
kUwFxiGVyD/Y3vXLmGwC/UOg5hdwwhBaXgv1IAmGcH1aaub+FrzepTaQ1vg3d6wb2M8vr0lWyN+i
n/JK15bE38a1rOdZE5hP7YUm1odCI9MC6blm+93w1c836PusibdcuP2m3euNbLFJ43yC0ghyYbZ5
ZuDdYgro5MYepsULMsmBpjthaGRbMqpEw5Ovvmwljw==
`pragma protect end_protected

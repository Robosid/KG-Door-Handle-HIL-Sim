// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yFFk6igDv5cr7piCJxf8HO7hYEqZExVAuJ7wW1yfxbb4Amo7QbznxIBUMK0d8qaw
rvIoQ5vBd6w7ZTe6O+WTPuHaTS/ayzzTqZU7C1KKGVNlCEs5horoVKjOHQdz6w9s
ckPxzh3/q3LSrBZrBA2eIA7yzcveBrSeEjc+C8Mrfh9UMQBz7cEf/g==
//pragma protect end_key_block
//pragma protect digest_block
TS4QFfK12bUoSsPB6UK+RphtwiE=
//pragma protect end_digest_block
//pragma protect data_block
wHDUzQbnfXhql5j/1cozW1qXCAyxMmdtOR7az93GdTczVLUIuE1Vr8oeb7yp0XYK
d2PCKlGLJ9Z0I9TGMGypCJNsutsQFlKU1r4YWcHLsMMAoPcdsIpuSK0la2NUkGRJ
FCs+ywuXZsYLYAtnrqHtdZaICgRBY5kxd8miNUNDUsSkuKHY5u1xMeNr5qpGjwry
W0VDA+O8Y1GyC3EMMpJBI0+xQqEmL5plGCosf0x55gzXFEQ8kfr84huOy8v0Rbx1
QVq7S4seZIo8Q4SpV0111VTG/J+l9DDaBbXl1GjfY5ammx60uqsJEaO3bnewquWd
dNtF0thk8ZNBsV6cUnw4qE0Bn258bcxQHgpOWI8a6Nh6mig5N14uyC3+WwPY6OpK
J1gwWJdvbeqO5W5ByuFb3Z1Gfk7ccKoBGm/Ed+nvHQSx75wDY/uF9ZrFb5YsXWrC
dGyTGZFISXTZnwzwxc5n1fDirkWgBuN/ZH6QmPsOdzIhVKaWyHiUB1ZUWdyyBLil
4+x/nJt7thY4bepf03pDMj/JNzPoRPEBmP2JIQooodiBacQvb7qERKEtWl/ycxMb
oyk8+fhQb7EBJptmOci5fRlskCJZUcqS+qJJuh7q4TtUNkKbk6znolNGHxmyFI00
JyIznjm47Y8s9VHl1DGTvoo0MZcxaMbmKZxrhoxVp0fWO9SIg1QSyKZG+6vgU2m7
AMro5sjjJiXUAM8mtPD5oICD0VVCiNPlF1CBv7/c+/zhtxaOoOT0ADZlzE0ZOAmf
fVrhYDxKvzsj+GykRsmApVuB/Kw/WrAV7hK+Wrwns8IyUman78AAoIeCoLCUcEQz
wNRoxHnEyd/aYttn+GdRTfY5PcZog+9z9ul0hV2eu8evLFT0Wn9rYWk4DJfXIxXP
WDiMjlgyjzIknZn4or+AHnt4UyeVtiWFTa4w9EaSJUc8zWnk1AN+xlPcUhArSwsY
TtLn1AMJypoCBPl0FuXBcz5NUJdV2YasDQF/GS4xDeDZG/pvdFqVO7D3Z5dog2jV
DgQa7vYqcBZSArFWrDX0LJT1kdsJFzprZhRqTF9Q51TM8eFi5gReYOOr/YqEd7SZ
ErnSznkZQtNOrfOrXJyxzXdMXifTYTNqBoPqOAOk5+lxmbEa8Djg/sfzB9iJtyAV
Ru70ISQEAS9AUeEBxCUkD47Dzen2L+asYyPb1vmYv1a3JPvct6rKsWF5Ptv+3pL9
GUN/70TOx3ZUq8SbG/rkgehex6DfAazzyTCwbaXIwcYG+RqeZRSM1+7Ofb7HadD6
Glds+I5crAME/njlVhp9HfKadUdMYUntQYZKSuWK6f5qzftsPz/iMWhFweQOa+6d
DHThiJ7WzhOCbVVlrQP9ECbLPTUwW+FwDDg6cp7h06wCy091PN9iHgpnefyMrJ3s
3tx1XtZ/OOGwkfqYaPhwXTPIIXLJGXUCVf/TUwJTGHHkNeaVc8ss6aA81tP4028i
jOOJWUXN242y8xWmJQHhTgupNIvhaa+E4wBdyY5EO+I56IsNMeRYWPHk0ndoAc2a
g0Qceooe/1slcuFLKQCGZ4Rmx256llO1wZAIXGGLKwPxa+7Y9zZkqp0ro/SkMiYu
UrbhsWfZcdHrDQRHOz3YRWF4TzVQD6TvZdrdm302LgBilOwhFeUDQW+5voCIB8xU
zzsCRHwSbBRHbv+ByJAir/FoJQSffmKVILivuHM6LNCnTPxn3pjGG3Ld7dWXmji1
8T2XoOACROAKn6N+/ivGWpXwfKg7zbCSwb8YUtXqikRzh5ZZsWggjlw3GaV8nha0
fgDAZ0A+23Hr2Sy7V3YWu4oOozjaBOELdRqapd1JbFdVCBBE2R35Q2iOOTOFQngA
wpSQwW9AG4PHfNR7BqxFdUUaAc0ttHMZ5CqEzgSD33Bw+9SnYQjIPkqyv+w5A2M5
BMy1E6nRn1y03YjJSyfE04/H2zO38vaVukqmXPnpckIdKf0KuppbdBT8cgksNZvs
th3cKktf86LR4F48oZCIfFZ46Bu+eB8FxqDJn5qa0OYD/5/rTnozbf67Q6EzzIf7
QGy0cLX3h9yNhcAdYyQV2MOj1KtvExw8ndbmGfjVayLek6X+rC8RY5Nq2bJbvlPO
OspA+/Mxp+iNdAVuEbkRf0gh8et1rA5UZoHwFzNbSGQcYiLstVVne4z/bDAtgWiV
VhwPwLTkc2fVa82V64zukO9CQliGmXCNlQZIshns623oIux87yrBqmuMXYTjLyU/
bOVlSrRn5jytFXi9po7IadgP5ovdcEZ07wUcNFMiMOAqZIiJEfd/VBBDP0vXk8pa
Ns3olR/Y+Iyrkh+hnIvNCm5HlJ5ZXkk7IMwRxO4se38qwKL4KHC0hzAgkQmbmsP2
/QbB5h2qusZRL2EQgkQ1lbFK1DnqFPcajsP9oKxKaXh/OydcnZ3XXa4OGynwyjUi
+ZfMNtASzK29ig30IFRSLyTH2E0cZIFyKN2D/TnDxqiTam6Ij4yct/UT5zwhXmG2
0jmMMoWyglOiu+4S/DC+F7Cnck7iu/ztYPoUNWi3THov1RwFaBrhYsOZkF5BkSYu
H8+f8MBns0wrbwC3/rb6/naS9bBgLrBQfjsRczszaqJkU7xuiCSuBSG3q/8jiD7B
SZfbTNLBO7rV25hz5cgvKHhhkWU0a3ZX/oawaY2+MvvKx0l3SIiJYAUrEwMy/3eF
1znjPzsHJKJi3V7HdQsZjfNnTHdwUUWeWQJAwvoLrmfL7sD2qhSqoY9l7EI5zWO9
fpkaRpu5lzATxm/itTBKpo7uc89DhJ8E2rD+An6NIjmyrvx1uXTzdC0h5eJPV0ip
TW13m8pXHi2CYIr0WvYVblT6Rkrf1V+ATKTFWoy9BxxY+OtwGgpeTFx3gzuINuHG
YJtq9frOydmxMkFM+86uH3ViKvp3BKMW53u+MXtfnvIMF6KKBoAg1Wk11qShNUA9
usxfV/Q1/hdwGsezxba4qHfoby1AnJn0+qvEHleKlIrmBYf3Rqc580R86/lyFwju
olXPEMIk33JYbm/hQeAEqpHvXg/OuvIpOgAChjv/20tAr5fdcOSzRmFrFDgubjNj
gLd9Au1UNIXmxBxFdLl6Zg2QgFqXNRBh/SBsp+yTVQmiAMUfYQkSD+jscR8XVq5k
iLWWENLsMO1Ggh5LlHb3QeO2/hj5cOD9vhGSU1ak8TnHdJnRBu4puWgAa4d6btsA
CdqjcJGiyKK1rF0woA6oUJ3oZUDVAruFEnWDSt6haCZs6g2ni3IimYxobqBivNG7
FUHiyv9Y1EpmzJ0OnhpSile86Atn6TMNea0AGULE0Ul3FkGSsAabKkcsfDQA2d/X
74RMz/GKxDIpWgWBrwnmy/Jfd9Wck2qDuZ1br1iXLDGMvqqF6x//xcrwaIcB2rpR
JuIo0p/pPGIpk3cehAvkOgmbnRMtKEqWlV/ID5Ohz6B6jtYCtyFnnA7+GxZBCalC
38aEKucTNjBxehK8sdsH7sH6iuRZ0e8jFMD0HXp4T99TmUb6hqmgJgDN0ZB0z9Xn
XhulLdNKg2GlPWgYg1VdyyKMpg7viRfCMhbG+W9YvQ/Mgt9bcNFXORbvh2NfnaM4
K7uRizWzisHphCDojWAjyFM8sJ98Y1ETsiKXiU1hiLmRgIQZPgaHIgkv7BqUJ9U9
mmrw6gpo/H8C0avlpGGwXA9pE8vy7OL0pSPmeMwJfxlq6gYQNDnEZthgOwvVfcnb
A97wWVihtGXKRywJgMPtco73xmI5KzYqQ4e+ZXYVAWfIVDcSlKusTffRGWTrhcmE
ZTFtYAhIaehnL2qUD5/PpjmPk0W/8aetfyi6QfOzRIpQ2dzV+LCSeJgbUnVuROGk
JTmbR/cfTOV9LzdOTobs9/35++g6c4NdN/daqwgvVPAtg60/7wulP9wi9VYFqFJb
m1OEqsBfMOOhwD/L4oyaH6FHeUM8Da7vGZbfIVKpIXVoZf07XpwoPXcs1BDI/0AW
EeqFFLlpebQ3cLW2KsrvD4Q1oZVZpj6qT8cui9K7drYLNBFxlk08ye9EhGVjq3xM
QGfE7sIZqxVpq+tf+zuMR5BnvTC6u5ewVk0+bdR7AnSUH6D8L5IxoOvA1Eh93jWE
BdDguoiZgWJzg0m599NYPp+6DKZLMGIea/BEMcgzt+zlkG/hptCxDNICgdrFlO80
NSlbEsZoFLv7/frLWwkq231Fmx9r7qY5ToF/rPq43xobTnI0MQOO74Z+ZSrMO30a
d0ECobCG8iLukFf+fECU+qLv+NKC4VB6sZDNcCvbM03mnDNVF2KC6v5HNy/zUY+b
Axu8F+akWMy+lA9+ygMNqTsM5Sc4TUzEnA0r1jdNxQV6CIPTKItsC3zc2/b6Zzf7
h/S/B7ZUvsfDo1eOFV7vhASex75JLK/58S4LJ5YGvBrIydFx+R27v5VWAVWUQTkT
8+uESopkJw47D8LNkswahKlI+daTzIt/bc8dm0GH1j99WT6kmSDMMSETedGszDaU
JUbgXopu31hDPBN+MJDNuGhtDbeIk1wejGxBHim9+X8pyeWniwKXc+rjYhGbRbaL
Qw8ptEahn3Q18CRdV/TFy6j9CA/Hw96QmCQa7ASdHtrGs5wTYlib6s+KQ/Kq4+Ai
d41/MgaamEWEbmcMuinZ3yQrqQ2GnwJs5xkZz93Drn3YDlIuwCMkxFVvtqW8QxlQ
72UGOBFbKoSyWz3eNj/4HxhYKwv/NI29nKgN++a8K5zR65dS/a2THvy1A/vgXT0H
EwHnjZUqRK6cJujo2n3Imy/9dlq6+b8LkXzL9r71CbaAya1f3moLtW6AWiZd2lT1
OhpMdxlX6nWApO1Z5Dmf3eLMR4LXkDldC+i9RcUs7uhf4MlXDeCcAgq3M9LCOAG0
Lb9bHm6shmK+WVhJ/ROe7wqESIrFy8bahPj73z1RrZR2YHfDGKLU8dcoP6OQ56ms
40JQDgX04wi/tSPDg+Tz7XSNjQEYMTCB+C+/AvlwySfq4Oho6p8x/8POkOVY9WBg
z31fM9i8ggZmBt7eu2/EWAZoI/rZ6WXKLVFtBY8ovtyJvL4DaAwtnT6fA2DBQinJ
oSvYD47qKRMA4sv6gsT41hxte739GCryhucEGer9VvrtDJkCvK4fZYgN459HVvKf
aOzyGGUGyaG4Yca7cLe9yjDCMWjLJ3WmWqfc2pI47oxHb4eK2CJg8Q8Q1ZVVQ5NR
VlGDGC3iK1wTh8B1xrQfjZAhocNw6H9R0twpXSZRvQ86wIVTSADoJdv4TlSY4fn0
qqWusbhhi4HVEAjT+eHEgMKiJ5rTDGzuB8ImqnQOnxj9xsUqga6LRsZyeVFM+5L4
myvx/8cUFtOqsDrHPSNB+NQi0c76qU/+tx4mO/goHCZEvMlJlxsc5qSicZVp8Jcj
ijP6C4iZeu3lW8hTqdJP+hXfBxjLPRejWWB6xJj6laBdMghh0yenXGU+9N3Rmsj8
la7NeYvn5M9GbfHD2g25urgWlCS87wDb7r4xwEqXLmnLT+RtBr9267mWmrU5eyeF
8NdyZK8S5I4xzNqKPDEO/+fpagIxJ5m+V65Sz+uqbNBwWUdob5u3HjqJwH4IxnsQ
vLxAc3FTPDtOpjh3r7ueTvPwXIFD9DT8l04jbT/17s8SVQJ+DCLw1AD+yQvlcK4Q
7ZMOqf2aHET5TS5d5/YrfPwGSEIeoqirGdIl2bnufRHwlDyYnzS1KYxniH1BYZnW
HuexDm3YxSsnDzzXcH8ZZ1ZeBGfaE+r8Bsmvp7nJN/4mJIA4pxVBaNUEG5wjgtel
+Zq7l8XCZq8Mna4GDyI1aN5yAwNIh+VoFjpgR8toREchaf0Z5zqeA27T7VThf77K
vT3NR6kcYC7OUh59RtrNVzhpaxQRihuh/AHPrKwP8APYWS7uRRI32CoItTWm0gmI
GuoXw5lXH57p/8B3zIH04Ee2AREAhYFshZeSIHsxWtLadTf4J7dMX/Fml5JNSMGT
8WuY/0R6Y7TtDeGuiApeH7NbGBzhPjqMoZvNDTB7ZewOoqfntTSm01zZK0sWXOeC
98VrN9aj//dxBnmi7pAgY8/lpQG8uIhr8+JbQSgw/6jBImvJIVTrGoiH3r08S0fr
YCZJifwXAvVzmWFDi4wB9UAFvPTwdGICefztyauou5fBxW7REr8wPi9nOjUe0e9K
c7qx+5+ocyzCNBkLcVf9HyUBQy16kqUBT7AIcPdg1A7LsHvznwzpkr5bQgVsxlm0
8+qWgauY2DtJtpuBriWumyiz1QQ8tTRGinX3dcGb9yzXqYGNsD35jVISZAm9sVqd
Cd/BuMmNrQrl/rbopTblNG3I/bs3iMi0LtL114o64OX4TeAlXK1Pu4rLdNd38Glv
zMha6Oq4noeqkQQ14S8JSJKS+2bVaerJ82LW6OpdPD1Kbkq/Szmy1v/WmzIhNwyB
2FGVqjEw6Xkj2lE7R39jWe/x7MIiKufh06RifbtLnYZiw6P9xg743ZJ+T5kgHyir
V8XTzBsYOdHDGSW4zYhWnCqDKi9Mm/PX/J0gOOLmYEap3yZg75mnBJrPAH6/tAnB
AGbDDDubnYYFImNS69GJyQFoyP+26JZp9RXtLu0GDVo0l7xGI+bNLmRiEQ0uHAZ2
bx+erOd4roY0kT2UUQ7C2PxkiFhXq7XZRN5PIUGLOEnnRjAinb1c8BOPWxpQCoer
4TQ9CMa5Pq2t9qEcafjZTmffRdbPEMMWkzdRLN19SUpC1LoZrL8hABDPs6fWK6Q0
YjTWXVuSgXerLhmjsjlQYzlPHfPp9JGW9MG1BdSHcrL50VK4CTMwm1cXHgtG1ZCa
x7ZaDPDKty9/E8b2bNAvd1AdKxFielfkXufK+crwaamnel6CO5nh5TsfAnFISewP
1mPlJJ4zprABeW4wrb55lvG1jwevCzM+KFDQKkwAQ2/0reh+WgDhgzhOZiaQowUL
mCfjaFZvEtYUoW8mEOloJkr/9fC6iQbLvGcl2jco98woXCGHudys1eJVylZikl8S
b/BYOeTctX+DUYOAU6yrYMseGRPLt4rYRcu8BNClTMah6BTxaqBra2CgxcORF1Mb
O3yZZHX8Hgl+caMrBrpYsoaZnQFFi09ycLxlkUWOzSUAStxY4QLB8dYqRcLiwYag

//pragma protect end_data_block
//pragma protect digest_block
IpeObODQ32Sux4ATC9g3/uTcSSY=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yAMIfKBlwAZdGKHHX5tp87SzkZy6VC+mB4dEXL9tEX8HBKWRW42JFRRvV2qeo83E
sRO4BsPEP6mGFU7wP0EYdZdTgq6ogxzUkiP9yJ4cAiCjzCy+WeJLcKZjp0H8aTY3
tIqcvmEYpPc47kr6eE/jx8PaPJ7j2uL18ySb4dC5XJXAcADSH2CBlQ==
//pragma protect end_key_block
//pragma protect digest_block
fo9Lbl4nNQqBn+sJYR6jHt8Ml0w=
//pragma protect end_digest_block
//pragma protect data_block
AVPVJrVgLKiUmN4+GcBvcGX/Lf3LrPGzLNsbbmoJibB/KjkbfsH+Gz2uKv88p8rU
d9viPBYkgziYhTOcOVjcillKyHdpL3FHxq1PPdGuGJ25dRcRP4cSm2t0SRYOKdxp
oHS9RxlijIqR5i6tYjyZBcrqwYF+sEwFbH6hDI+K5q8cint4ARBVKWAxva6kfDSP
fknmfG7GVk/3cIAAuU01hh0eGEUqOrif2HQn2TQiL+bIl42ixoJbNFw0YzNy2t5E
2xDrnLg29avax22CXmfXjgOEfVhRohbOuk8Lrv7YZ+NkFTBDAs6gnJhEdIVMyttA
Gnf/ElLR/HbRdKO8eMgCjtGmR8AbZqgQ/mQHVkRJhFIktrua3WsTWaKbS/uS4Zrd
Bt814YMvl0RSngyJw7dPm3zGq/KKrvO3GIIS48QZ2IyeabULMpUjhfVBIAkvFVEP
Rkf9KDsEr7jPXEWOGFmeve8TVAXqN8rooRyjJpuDNni156v+LfQVYs7z9tBu+20K
3pQMkngaWZhYRKt5cRwJ9maJLCKmtKEzfmtsey42iWOk3maSpWjg1A+w9jl32qpU
/OvXt01yNXy1y7la2aebFA/hz8C+zIy+VCuHdvrSWIeteyGOVFvE3gc0NDmBPo+5
BXAgyXFnPFovwpG9BJ3qDG7cdqd4lgNaM7J8dCMndMz6FNytuvcboyrijtvtbigz
a2gm6ALvAviIUZLDfKsurpxRjqttxVNUm1cSKWVIwlrl0JFe7kdf2EDxaxjD8jQn
JicajSN14tfCyqxayogILS9DumWhyfPgvZbiC7JMTwrhMlCkbJCddfz333s5zMWi
U8cvBspDAEtvrJk23cjoSX+hvLBqhbi5ii2hWBE0yb2kRvpXOtg06g44W0znPp0M
euB96TksQ1Nslk8D5zC22KJz2GCbj2i5iQN1CIhz5YjPTgziwVQoFMit3q/Iv0yP
Pm1RzHRpPj00d6Z/rLT1To2hVhrAW1yspQkkinSfu5FvwVyKozw52swYea5WiRP5
7z2ny1DK/BcUmL5rm4AJvHUX+6rK81PMh4fWlNp3oE3LoWlACb4tmuiD+7OG3IpF
zQPy2IGtd6XFfnAtMI/UhShg4RU/Unlw14CEI2Y+0PINjFSofgbMEY4HWDSszRgy
O0FxBuwSfFLpRx1aZN6xC6zBfDuJQnfVlU3z/K1LzJ1QpTVaBdUnfS98XDIq8LiY
uL/laHYMjdpzM1kPdz3KUn4qUBvXA4JunUJStFoUjN1JSWFGdHdJooCu35JB09n5
UXHWNHZx1iMPrhkT3lILK5yPCF5yX6Bk9N0d6NhoPcq9AW2odQCOOnZMLfum9Mip
NvhcZ0pHlZ0eO9lRo+9gjoJJaafC1NV5PjtyjIxKw1edRcikdP9Jj8RenZ9SYX3g
+oyS3LhPS76dYKPMUHFllYVR+McfVhCPxF1dQO5OprKDhGXst6/9qHObqzGZsMLh
zZpWej6tsb60pF96qbiIEcTa76T53eqjESB5pF42BWMeMnqHbcPyX2HwJZp+9HxA
ObLTL0YBqHzanunsEr5DPA91tL2X35v45RaOBlFoX7gzLvCgFOdIbUPx7WZVdkI9
Fc6aH0erat3CWUa0Lr0rgxbtkhoeZ9hzcqQWl0Fz91Fmn2MkShxzevO0v0YT1f2p
JkECQbFQ3/TekDINk+VoqwxgQdipyrJF/15Fj5IXeES6IYfqlCEthwS5560pBAje
B9YApQjJT6bVEzzYmqlxEwDUgbaNNFXQW+d2H3+HLSbh557NYNv+yAp6kwHFR70j
yAec0bAtETcK7lAaruw5LkElj9TLKkQRoWt0ytakkXcSNxyKnuNGq4e7FekIwFOU
Bvi9R3nJCUg7K/MR6r1mC7s4sTeV2l/RdGuLgggscj6fRAuNIw+vXmlRruox8k+p
ECv2PD2S00Sw4Zn0OwaUE9kNHAqdH7YDEJnzSq9vIurBNkVDPh3rwlJgWZ2vNdzK
fhh9BhoiQp6K43MiX4STg4MV/SuIsKUQl1h/Sw1H8H5El+AqYa4FmVj/6MnUG+ga
H1flkbe0e8uslivsFa0fSWPkPJrbtwvWa/4E+OVsxBxqbd9p+ZDdHOB6qs7A76YM
efY4344zWghcIUCB59lRqjYmahS9aDg0jm0h5RIb9fX4e5MysVXIQLj6FOh5axxO
UTzlhYO1Z94h0GYENUNYuc3ZnRbjwHw11O3nemV1HnB7T0AABr0hoWrc+W+fn13U
ZC+th9PbNDgR1s6h2F/LBRvKCyAOI2PAmQZo0XHAzXWa/6/gXiX2W3as5w+nX+nV
GOdkseEezNThpqNFx+D6yxJ10v05Syw2zfhg0AdGM+Xu4x6k8b1qWvGLwWAmxXnT
fl/yKq0i2u9SzcPhM5oQcWPfq5r29wl52edXY1lvmtMM6g0bO6fKvF4eM88k0e8d
KjtUYBQusajDGnt1GMARcrAxk2ZvdLh3AZONodjOdxCWlLnYCq3QPnmoWFht+T+L
SfPfOSuxdS9/N2Ikkzz+sXjOKWAV5PZ/OrCBqyGmzPmdclqwiylc7Nx+Y8Qb5/Y3
sL+I32uSmnLo+f5HlLZ5geoaGL4RYmYIJJHRCDnKDgy/kpATw1WHElSc8TFL6cwT
MZe8E5+r+fe5Qh7LPXakfIVXAG/PpEyrMnT0YgeSAfwXieAYWG3bbo71Yn7oDR9I
+ZfcUfVrzrBs/ZDO1A6shOAwbBvgvzItsEZRc8TAHSugVKU4Dl21TJdatkVP72rd
rzqRyILsSiS85oRdivGR4AIDGPbftmwy2g4ovFrEl8ZtWn9c6KQG+MDUc7vd4FNR
BmgCLj2ROHGwmXqWM5jGHEa9aVIMdM2eqTxb9CQ+rMby3bgyMSbZfLbJSyeqUQa1
J6PJygzmI+qPM6+Pt8YVk6+Ks+Eime7kzUvLRuBlBypwQ2bG6oYt/kOBbx1jTsjX
EesV0UhP6aN5sDwENs4fP7qIpcNXXQvdSlkDVRes8gKSlDeZfg5CjdZhPfrwiETU
eUW7SCF81Hpqy47nntPAuYvwUmZ6sPZ7j75+8kBRX1JEYFvGhsmO1O6Y8Tc3BldN
VSwmZ5bvNmYX28SyJYwLIk/Iu/bnO+ulHE8Cbm+NnYoJAFKB5JChPGR84mABkrOa
RzgvccpiWr0qB+g1c6pskpqfpM317SVpKBqx60niEjrBdAu/KcnHVl28MwufqW2s
JyiWhYPA4YocZt3p866RKeN1eISjEvANxtS3jJ74+g/Rm/QSdKRNudPvYPO4VaZ7
2/yOwxx1A50TXodnNo7SgVLO3dm3plNeiIwUBgSK9wU1MG0IOj6jEEI09wZ4hQzb
C/qnJV3y/KA39M5LsCUqzLlWMokwm8YhP9j0gm2oc54rl0BsJXyCiKVyQS+NYOqj
MIgzddwOcmYrNLBPN6d/XmpddVtktLUpoYDEPaMai2fg/KsN4JdBAQCIQyB3+p0I
SiB0fSsQd2Cw1df109N4BHGuykP0z9ozQLkbeFykVw1BJ6O5TuVqrVeiRiCZJjxe
4lfigu6HMpxUlDNoLHfxWz0/CN8PeoXQY6OobPkB8FeNV6VgqP8keBCX0MzYxtgt
nUnbGvHLTwcgGKp6y6yQwbAlbg3YAtlCXoDv7Xy1BpjdnkbDjwoxIOYM9IWwMuV+
lVUZmVIbLotFvNTG883OzfvGsbVFOBW3RTLmMIJWez1fg86xPuu8vbMUCcZizOG/
9GOzUGE9mWOIBq7E8J0SIpE+gfbMlliWgiUnq1Kl7cVDYYebznJMK6eowbs6mSCE
8UOvkKLXzAWyOkSoOi2+lqGc9SiJWxeOmaaBGamcXyVQHmxj/OmcrkiElZshL5bJ
lhPgTJNqIiGPZMJAYsvLYMXzNAkNtLBWlxJZD0xVtqmdZZV3QMUf6sLsSykPOt2g
Vc0l2SNIi86Z8eZpFH7u7NQqD006akkiShOLrykykOz6Bzsfot799fwuponPfxPJ
FRrTp0ASYw3bLbLPnWuwoMZj2y1KE+yCklEPq760xjFv1KjyOXPDwh5AS3RlbVrS
Zyt7Nmj1ZO7U64IVQFryGsez1QSNlfYdzG7O64aiW7SGGqs0+hDXhnoXDTLVKw1s
6z/X0JM6XWoKMyXNQjeC+yUZAAQ8tT6MutMSIWTeulD1KSbTKd6eTvGt7+sprawh
zcEBfkIxDgn639BdSoiNHVy9Uw96ennh2bhgxG2p7hbwIE06cOFT/Op9APC5Jcsq
ju9nXoYRiep5xqbXYTfVCDRuC2nKhLt4oBJHtUixN7XJs4WsIFzpWaoaUH5RkAc4
3ImWpcLZAJodaqJnuC1fyjSHWUH3s0bwnh/Ao00JjpPEbF+q6qFURgJN5K4RHu+4
21zKHl30NPT6moqgkqtMho0jMQcpjJ5+m+NOdMpffPYWFocs4xSJLvwLtPk0cXUr
qmrhzK5F8NBiNK5HBi8qL4dNH19alsCZkgafKXzxm/Ly50fjWmZ5iMKZk+DZ5Zmc
s1HsWRW2N8RC8L3SV6lMNyRnJHJEBjigKC4vi7gAUoHpPpvXmX7qVy0Kl/TvKNVA
BGYHPTEZPFRkitL4fTkEXqQncG/eOlVGgM2Ex5Rsw+BuuhOTweUBOffIcSCcFjkH
CjrY9C3cEjKqHp+GC/Vh90uU3WuICocqMJn6oFN7qo3KUo+hew9G1/cxUncQuUG4
ti6C4m+yZux9d4J9KVifQBHxMXSVx/biEhzjvW6FUhmdSOQTukZQXfMdOd+kde7q
+o9l/eIFcAw3i6etyvD0jaHeYbDG/tf5NwRA6DdP7monO2kxGkazwAOwFlEajhyW
qkWk7NzpGVseHkpkYESS0ndWzG/II4zMAzwJKqJ4GKkglxqzSdoirR/joXVFKOBk
mGwPseZg0QYC1blkTqYcMfdtGO/ar0QM96rTS2OP3mLRPskWRum+N2OsYnbMtZI0
te4selrETcwGDtcuT0F0WGjBaig+Mvt2HcEhULltYFtspqOZlYwc8swtPSbqStiU
Gu71QG0eBg5ICF+FU0nab7yBxcsrZ8wXuO22U5EDtpFCEqBMYfOiAvU/zJNabCWz
+k5ROqamjpqTxS8LH7/MzC9zBzae6+phGLb6esLWvHBi1ZCjwwyMKiio9zRd8n5D
8uGf6TE2dRtzRC8jGBLevPokcxDy+cvMSlN0YczcIAIoqhTFZpCoDxCoU4iPR6OU
Thh63BicKB/XFHMuF4GO/psnzFMgfM2IUiVTCU9UDU0XZcGzy9eip28Zrcti52po
oUQom5SR/SoYmFe1W7duIWrJkdlQuAYO67ObZHwGDonDtoCaXM1pkPBgjyzyoqW/
edCgssslbKU9UTB8CJSqAHgH4R8GGE11QWC0qGEfVe3En23ci2ZZbGl8uBjYPrvn
V1A0bHWP/L/pgyuTq/3xUw2o/LnbAT9ZEOqmUpbH1fY6/vt64prQ7o190j0erPQB
NPRJW8g/jCkn9ZPB9LunZu0YNRN6Nk31dU2RYZQonLMgkIRWvb1L3Llunupwuwaz
W84K0/jYv/19GPr6azpt1TOeiuMGPNcKD5sJIdbmAcEjb7Hf3A4bX57RC43esbhN
rs9+XH2u4mBRXU0l4bkTOMk0JwUpDyJrsBQwrB1Ap6EQ6GYh1cQni2J1y2uDqNBg
1TUz8TKf0S4r0yU2WH+IinO4FcEjmjmFN4cE7pF2pVBPJIPoaSWA7TxE2WcXh0WJ
ElIctP/b7BOV3UYX3mP4t7MlBncRucFQFlTMWQAUr0fJDIyD07cbdDD1DdZXBrbx
s5BSdB93WLAY2p4zYr6WnT3lU2JI7LUlp4LSOV9i4ER/iPdABjBpeX0FxUuVb+M9
2OTPXG1MZ07QH0aZX9gfOV3IrFokE/J3jd1zkJZNcF18R9bDQEJjgEmoECYS9bB5
uWCxHV6m85T6L2wrc/vQg8BMO+GJ5GNaWAKMumNmlr+DZgXqXOweoFFEbGu5N+SY
R8ZbhvPCMCzzoyzTo5yo9a2bEoU3y4Hq1AhInn17YmSXYVUo3HHmgO4Pbmw0Z0MV
i+LMNVyvtEZdipAWpzOeEY9DKEzOGia9lLSswj8S93taeY/cbRzQkZeqnTFp5LTv
bTXLFvtxJeY5bHWMLR2nWGWSJB9fATCtj/zCayZtZcnCy75OUmpef/wjOMivCdcW
Fo+dnPOSEdxvRsFEeRwDSwTA/RZL0s0AcYaB/F8LRfq61e3mtHB6Z2Sq23HGiTrk
xA2apxnG3jqwlfj/0qOmYK4K69V8kJytNiI0QV1xpNGdqadtigB8ENdHGrhAROoe
ziXVd/simdHFo6DZjaWMuLrcseHzZMEUbPzvFkiGyqytLC9zaJLOP9r0DjYgkffZ
AgOhDyawRM+Pre5ordN3vl2QqG2Vgtb5L1PQStUnoVy64DEnXFq5kLVMUgDxZ9mm
h1yNmQTb9vMJ5qkA0f0YsIFouprgUTBhC+Ed+2hzYMSmHYFw+H651QmFtbjVEyWZ
RJlf5zKN8B1w4TBpOjWiTEKykch6qggDQtl/eGPKVUI7FfBmgPzneB5RVVoEY518
fXm7z25MAdkyHL7RgPdSSTS/eWkcmRdB7brlmc3ydsbFNAg4zWikzRVx+oTEHUqA
+u/O7+lWQ4VTo9FAYKu85KS7LYRaeFcFcGQ8QxGhJSW3Z7yftToSBtbJccx7psJP
qa3Fh+gI93+hLSS6hwWWtlaztlA9Ds1689x+kDPgJA/A3nu87LFnkYQAQf8zRQ91
gLlcWDDaZUM8La7R9KUiMmv8clpZlT5KtXhr3wEk7DXfzrD5QaUwQKdbGU7B6jKF
6EnfY3hkBXp9rC88SdFwrGnFYIpSw0wIt8CRnNik1RQF8SE0QqemMPpfs2cexyKr
6UWHw97xwkme+gVaJOYh514Qpi1mm0bewh4wtyG++Z5KdftlMCRLOkyF0ImwEr+s
L2ipqEkn8tVPKpaMe1Y6k0K6zyBSUjkut3mhopNGQOEbbE5dsN9SP24wlErMqjjp
J8/aLjgBemwpSFt2RLN/UNS4bcePh8XPG2j8ozYIocYV1IhEM6Oe4aHXpREGzu3d
RQxGEGLCbNKeB+Gcl3IYwWd8Wvo0ZQ8aojftAX7hGB/sS4PQ+mINFJsb8WtZ7z0Z
CwkufkftNgdIS6K34V21EcKMPbWSO4ShX4W4V2gXd9xnqGtGW28U53Ee6wMdCycB
95M+0P6OOIU9ah1XDW79XGUgYnMa3FzipzVepFevPmu0z8SXRs2QvY6mAdSudCT8
ppL32+1I7GLSxQw3vYbsXpE8GZT/yA7Zj3EJ7/0GN9S2aw21P4mDT8AwiCJnc7Gp
fba4WEwoHDc6+fsrTu/U198SSjnE+mpAMgIHX4qq2kvxNb/HVfquFYETCblMv9i1
ai94faP+Fc/CwN3Wq6wCx//L0meddP+WEMz0G7183A6Mw+NN8KkVoCPJBS/iH306
nMcunlfTdmSv4qPksasuUibVtNTeHQvTlWaoRRvcTNKU5qZyzlFHzZ/IeylV36id
GgYmNxpVYUhOPlKdDCVTgkqMnZyQxr1Vaxuu9Y2YkRa/009a+7VNHsq4UsX2rR45
QdYK0et+czvlGWyQva6AFJWn3PRS+IK7OCwFCZRaCvLMPuYYFaOAxXkA/JvUe5E+
Tq5b7l+gi1oDEBy7u9QOctyhtImlSXmsqg6H+5kAyWI2MXPX1fUXtcPJ/4qs4YbA
vn5GRRRBjtM19D+PAZSyrTSuM1x6RTgVzueUFxp+39UGfLgbmhs5HXSgodZOkObS
7oUujBjaeDXVbnP3LwEZ0LhVUy6anLmdg1e7zctAei12BAcqGhP8hUXfG3CoOAyS
XVO+IazdhvyDDjUuuhBLDj82GNMUDsWG/1vCEdozkI5pigwx4QZ0Ypb/ncieDBc/
snreU9OG0hZOOaoo4d3cNvN1PUVdeF+ljApSpmLIpUGfHOqJ6waRl3tF4qxgTQHM
LfvB96k1dHThM3Qb5geRmbT3UHZQzVmYCdZVCQGHA64bicAxG024zVvuekFwAosR
Wf+PIutrKPFq1BOd1ul0Vbzqzkgj1AUQuxmYszziNoAppVONsRAeaoWPYQ7c0Kkl
owKNxf15CV3tIU8TLlJF1cPDl+oLCsBcvLkIOfoCAj5JXCVMWfFH6HaY8r0UScs2
tqSULgkNchGeAp0pJvP0+UhdH2BbRoaphx2urFm+32/47kcAGtMXPirGAcL2i5kT
XtM4WRcmwEg2cXdM2JRE3YNL20eSC8EzEoaTDazIIxQrm4ud4/bLNRvvEXuUrnui
BuDKzdxa3mfEMGQcqY2Vgzjha09egpqt+vK5s8OJ4uGF4Zrc4Ygy/MlWL1CFBXlM
vds9BRm3TPHwJAfa98B0zxFYe1T6qe3kIv+GdzkhnyGIEiDFTlEfjTl2tPe2u8VR
AtFmcEhhFYUXXCJ7sjNh9G8jImi40dXVLd/SuRBsHFf2OER05V9VR8uOMIKIsStr
pXHwVW0YpbK+LinoAZCo8zCJhzh2xqvcmAfK6pGMGit27ySLmhg+R1wKAz28/e4E
SQGfXHWI03O6IAG5fUFcDuZGWZ+0kFULoqEc4i00gVZy+LGpsrj+Yo0TcXLTi8o0
YoWus/lf375jrW9jEE6a683e8Gm/WlTFVey/MEJ827Vc3YptdsKrlEYkZnIICin/
D1shr3eX4NiGAlskWLQGnN/Q7qOWvKyK2Xtlwzjf/OFfcCwkaJFi0qlj9VSLQyuN
x3gxcMZK4WBxVObxrfuOdoGG7ubBd4QchnYl4w4Qh4vVhh5qxI3D7h1pf7omIzNR
oy0t7SpTTLrTkN5otAFp/P6vaCr2BgyoAsR5xnpy+mU=
//pragma protect end_data_block
//pragma protect digest_block
HCN3GqNya2Ul5uIWB9nUlQ/M/M8=
//pragma protect end_digest_block
//pragma protect end_protected
